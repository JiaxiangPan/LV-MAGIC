// Benchmark "top" written by ABC on Tue Nov 12 20:13:02 2024

module top ( 
    \a[0] , \a[1] , \a[2] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] ,
    \a[9] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] , \a[16] ,
    \a[17] , \a[18] , \a[19] , \a[20] , \a[21] , \a[22] , \a[23] , \a[24] ,
    \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[30] , \a[31] , \a[32] ,
    \a[33] , \a[34] , \a[35] , \a[36] , \a[37] , \a[38] , \a[39] , \a[40] ,
    \a[41] , \a[42] , \a[43] , \a[44] , \a[45] , \a[46] , \a[47] , \a[48] ,
    \a[49] , \a[50] , \a[51] , \a[52] , \a[53] , \a[54] , \a[55] , \a[56] ,
    \a[57] , \a[58] , \a[59] , \a[60] , \a[61] , \a[62] , \a[63] ,
    \asquared[0] , \asquared[1] , \asquared[2] , \asquared[3] ,
    \asquared[4] , \asquared[5] , \asquared[6] , \asquared[7] ,
    \asquared[8] , \asquared[9] , \asquared[10] , \asquared[11] ,
    \asquared[12] , \asquared[13] , \asquared[14] , \asquared[15] ,
    \asquared[16] , \asquared[17] , \asquared[18] , \asquared[19] ,
    \asquared[20] , \asquared[21] , \asquared[22] , \asquared[23] ,
    \asquared[24] , \asquared[25] , \asquared[26] , \asquared[27] ,
    \asquared[28] , \asquared[29] , \asquared[30] , \asquared[31] ,
    \asquared[32] , \asquared[33] , \asquared[34] , \asquared[35] ,
    \asquared[36] , \asquared[37] , \asquared[38] , \asquared[39] ,
    \asquared[40] , \asquared[41] , \asquared[42] , \asquared[43] ,
    \asquared[44] , \asquared[45] , \asquared[46] , \asquared[47] ,
    \asquared[48] , \asquared[49] , \asquared[50] , \asquared[51] ,
    \asquared[52] , \asquared[53] , \asquared[54] , \asquared[55] ,
    \asquared[56] , \asquared[57] , \asquared[58] , \asquared[59] ,
    \asquared[60] , \asquared[61] , \asquared[62] , \asquared[63] ,
    \asquared[64] , \asquared[65] , \asquared[66] , \asquared[67] ,
    \asquared[68] , \asquared[69] , \asquared[70] , \asquared[71] ,
    \asquared[72] , \asquared[73] , \asquared[74] , \asquared[75] ,
    \asquared[76] , \asquared[77] , \asquared[78] , \asquared[79] ,
    \asquared[80] , \asquared[81] , \asquared[82] , \asquared[83] ,
    \asquared[84] , \asquared[85] , \asquared[86] , \asquared[87] ,
    \asquared[88] , \asquared[89] , \asquared[90] , \asquared[91] ,
    \asquared[92] , \asquared[93] , \asquared[94] , \asquared[95] ,
    \asquared[96] , \asquared[97] , \asquared[98] , \asquared[99] ,
    \asquared[100] , \asquared[101] , \asquared[102] , \asquared[103] ,
    \asquared[104] , \asquared[105] , \asquared[106] , \asquared[107] ,
    \asquared[108] , \asquared[109] , \asquared[110] , \asquared[111] ,
    \asquared[112] , \asquared[113] , \asquared[114] , \asquared[115] ,
    \asquared[116] , \asquared[117] , \asquared[118] , \asquared[119] ,
    \asquared[120] , \asquared[121] , \asquared[122] , \asquared[123] ,
    \asquared[124] , \asquared[125] , \asquared[126] , \asquared[127]   );
  input  \a[0] , \a[1] , \a[2] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] ,
    \a[8] , \a[9] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] ,
    \a[16] , \a[17] , \a[18] , \a[19] , \a[20] , \a[21] , \a[22] , \a[23] ,
    \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[30] , \a[31] ,
    \a[32] , \a[33] , \a[34] , \a[35] , \a[36] , \a[37] , \a[38] , \a[39] ,
    \a[40] , \a[41] , \a[42] , \a[43] , \a[44] , \a[45] , \a[46] , \a[47] ,
    \a[48] , \a[49] , \a[50] , \a[51] , \a[52] , \a[53] , \a[54] , \a[55] ,
    \a[56] , \a[57] , \a[58] , \a[59] , \a[60] , \a[61] , \a[62] , \a[63] ;
  output \asquared[0] , \asquared[1] , \asquared[2] , \asquared[3] ,
    \asquared[4] , \asquared[5] , \asquared[6] , \asquared[7] ,
    \asquared[8] , \asquared[9] , \asquared[10] , \asquared[11] ,
    \asquared[12] , \asquared[13] , \asquared[14] , \asquared[15] ,
    \asquared[16] , \asquared[17] , \asquared[18] , \asquared[19] ,
    \asquared[20] , \asquared[21] , \asquared[22] , \asquared[23] ,
    \asquared[24] , \asquared[25] , \asquared[26] , \asquared[27] ,
    \asquared[28] , \asquared[29] , \asquared[30] , \asquared[31] ,
    \asquared[32] , \asquared[33] , \asquared[34] , \asquared[35] ,
    \asquared[36] , \asquared[37] , \asquared[38] , \asquared[39] ,
    \asquared[40] , \asquared[41] , \asquared[42] , \asquared[43] ,
    \asquared[44] , \asquared[45] , \asquared[46] , \asquared[47] ,
    \asquared[48] , \asquared[49] , \asquared[50] , \asquared[51] ,
    \asquared[52] , \asquared[53] , \asquared[54] , \asquared[55] ,
    \asquared[56] , \asquared[57] , \asquared[58] , \asquared[59] ,
    \asquared[60] , \asquared[61] , \asquared[62] , \asquared[63] ,
    \asquared[64] , \asquared[65] , \asquared[66] , \asquared[67] ,
    \asquared[68] , \asquared[69] , \asquared[70] , \asquared[71] ,
    \asquared[72] , \asquared[73] , \asquared[74] , \asquared[75] ,
    \asquared[76] , \asquared[77] , \asquared[78] , \asquared[79] ,
    \asquared[80] , \asquared[81] , \asquared[82] , \asquared[83] ,
    \asquared[84] , \asquared[85] , \asquared[86] , \asquared[87] ,
    \asquared[88] , \asquared[89] , \asquared[90] , \asquared[91] ,
    \asquared[92] , \asquared[93] , \asquared[94] , \asquared[95] ,
    \asquared[96] , \asquared[97] , \asquared[98] , \asquared[99] ,
    \asquared[100] , \asquared[101] , \asquared[102] , \asquared[103] ,
    \asquared[104] , \asquared[105] , \asquared[106] , \asquared[107] ,
    \asquared[108] , \asquared[109] , \asquared[110] , \asquared[111] ,
    \asquared[112] , \asquared[113] , \asquared[114] , \asquared[115] ,
    \asquared[116] , \asquared[117] , \asquared[118] , \asquared[119] ,
    \asquared[120] , \asquared[121] , \asquared[122] , \asquared[123] ,
    \asquared[124] , \asquared[125] , \asquared[126] , \asquared[127] ;
  wire new_n194, new_n196, new_n197, new_n198, new_n199, new_n200, new_n201,
    new_n203, new_n204, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n211, new_n212, new_n213, new_n214, new_n215, new_n216, new_n217,
    new_n218, new_n219, new_n220, new_n221, new_n222, new_n223, new_n224,
    new_n225, new_n226, new_n227, new_n229, new_n230, new_n231, new_n232,
    new_n233, new_n234, new_n235, new_n236, new_n237, new_n238, new_n239,
    new_n240, new_n241, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n280, new_n281, new_n282, new_n283,
    new_n284, new_n285, new_n286, new_n287, new_n288, new_n289, new_n290,
    new_n291, new_n292, new_n293, new_n294, new_n295, new_n296, new_n297,
    new_n298, new_n299, new_n300, new_n301, new_n302, new_n303, new_n304,
    new_n305, new_n306, new_n307, new_n308, new_n309, new_n310, new_n311,
    new_n312, new_n313, new_n314, new_n315, new_n316, new_n317, new_n318,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n417, new_n418, new_n419,
    new_n420, new_n421, new_n422, new_n423, new_n424, new_n425, new_n426,
    new_n427, new_n428, new_n429, new_n430, new_n431, new_n432, new_n433,
    new_n434, new_n435, new_n436, new_n437, new_n438, new_n439, new_n440,
    new_n441, new_n442, new_n443, new_n444, new_n445, new_n446, new_n447,
    new_n448, new_n449, new_n450, new_n451, new_n452, new_n453, new_n454,
    new_n455, new_n456, new_n457, new_n458, new_n459, new_n460, new_n461,
    new_n462, new_n463, new_n464, new_n465, new_n466, new_n467, new_n469,
    new_n470, new_n471, new_n472, new_n473, new_n474, new_n475, new_n476,
    new_n477, new_n478, new_n479, new_n480, new_n481, new_n482, new_n483,
    new_n484, new_n485, new_n486, new_n487, new_n488, new_n489, new_n490,
    new_n491, new_n492, new_n493, new_n494, new_n495, new_n496, new_n497,
    new_n498, new_n499, new_n500, new_n501, new_n502, new_n503, new_n504,
    new_n505, new_n506, new_n507, new_n508, new_n509, new_n510, new_n511,
    new_n512, new_n513, new_n514, new_n515, new_n516, new_n517, new_n518,
    new_n519, new_n520, new_n521, new_n522, new_n523, new_n524, new_n525,
    new_n526, new_n527, new_n528, new_n529, new_n530, new_n531, new_n532,
    new_n533, new_n535, new_n536, new_n537, new_n538, new_n539, new_n540,
    new_n541, new_n542, new_n543, new_n544, new_n545, new_n546, new_n547,
    new_n548, new_n549, new_n550, new_n551, new_n552, new_n553, new_n554,
    new_n555, new_n556, new_n557, new_n558, new_n559, new_n560, new_n561,
    new_n562, new_n563, new_n564, new_n565, new_n566, new_n567, new_n568,
    new_n569, new_n570, new_n571, new_n572, new_n573, new_n574, new_n575,
    new_n576, new_n577, new_n578, new_n579, new_n580, new_n581, new_n582,
    new_n583, new_n584, new_n585, new_n586, new_n587, new_n588, new_n589,
    new_n590, new_n591, new_n592, new_n593, new_n594, new_n595, new_n596,
    new_n597, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n686, new_n687, new_n688, new_n689,
    new_n690, new_n691, new_n692, new_n693, new_n694, new_n695, new_n696,
    new_n697, new_n698, new_n699, new_n700, new_n701, new_n702, new_n703,
    new_n704, new_n705, new_n706, new_n707, new_n708, new_n709, new_n710,
    new_n711, new_n712, new_n713, new_n714, new_n715, new_n716, new_n717,
    new_n718, new_n719, new_n720, new_n721, new_n722, new_n723, new_n724,
    new_n725, new_n726, new_n727, new_n728, new_n729, new_n730, new_n731,
    new_n732, new_n733, new_n734, new_n735, new_n736, new_n737, new_n738,
    new_n739, new_n740, new_n741, new_n742, new_n743, new_n744, new_n745,
    new_n746, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n835, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1005, new_n1006,
    new_n1007, new_n1008, new_n1009, new_n1010, new_n1011, new_n1012,
    new_n1013, new_n1014, new_n1015, new_n1016, new_n1017, new_n1018,
    new_n1019, new_n1020, new_n1021, new_n1022, new_n1023, new_n1025,
    new_n1026, new_n1027, new_n1028, new_n1029, new_n1030, new_n1031,
    new_n1032, new_n1033, new_n1034, new_n1035, new_n1036, new_n1037,
    new_n1038, new_n1039, new_n1040, new_n1041, new_n1042, new_n1043,
    new_n1044, new_n1045, new_n1046, new_n1047, new_n1048, new_n1049,
    new_n1050, new_n1051, new_n1052, new_n1053, new_n1054, new_n1055,
    new_n1056, new_n1057, new_n1058, new_n1059, new_n1060, new_n1061,
    new_n1062, new_n1063, new_n1064, new_n1065, new_n1066, new_n1067,
    new_n1068, new_n1069, new_n1070, new_n1071, new_n1072, new_n1073,
    new_n1074, new_n1075, new_n1076, new_n1077, new_n1078, new_n1079,
    new_n1080, new_n1081, new_n1082, new_n1083, new_n1084, new_n1085,
    new_n1086, new_n1087, new_n1088, new_n1089, new_n1090, new_n1091,
    new_n1092, new_n1093, new_n1094, new_n1095, new_n1096, new_n1097,
    new_n1098, new_n1099, new_n1100, new_n1101, new_n1102, new_n1103,
    new_n1104, new_n1105, new_n1106, new_n1107, new_n1108, new_n1109,
    new_n1110, new_n1111, new_n1112, new_n1113, new_n1114, new_n1115,
    new_n1116, new_n1117, new_n1118, new_n1119, new_n1120, new_n1121,
    new_n1122, new_n1123, new_n1124, new_n1125, new_n1126, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1208, new_n1209, new_n1210, new_n1211, new_n1212,
    new_n1213, new_n1214, new_n1215, new_n1216, new_n1217, new_n1218,
    new_n1219, new_n1220, new_n1221, new_n1222, new_n1223, new_n1224,
    new_n1225, new_n1226, new_n1227, new_n1228, new_n1229, new_n1230,
    new_n1231, new_n1232, new_n1233, new_n1234, new_n1235, new_n1236,
    new_n1237, new_n1239, new_n1240, new_n1241, new_n1242, new_n1243,
    new_n1244, new_n1245, new_n1246, new_n1247, new_n1248, new_n1249,
    new_n1250, new_n1251, new_n1252, new_n1253, new_n1254, new_n1255,
    new_n1256, new_n1257, new_n1258, new_n1259, new_n1260, new_n1261,
    new_n1262, new_n1263, new_n1264, new_n1265, new_n1266, new_n1267,
    new_n1268, new_n1269, new_n1270, new_n1271, new_n1272, new_n1273,
    new_n1274, new_n1275, new_n1276, new_n1277, new_n1278, new_n1279,
    new_n1280, new_n1281, new_n1282, new_n1283, new_n1284, new_n1285,
    new_n1286, new_n1287, new_n1288, new_n1289, new_n1290, new_n1291,
    new_n1292, new_n1293, new_n1294, new_n1295, new_n1296, new_n1297,
    new_n1298, new_n1299, new_n1300, new_n1301, new_n1302, new_n1303,
    new_n1304, new_n1305, new_n1306, new_n1307, new_n1308, new_n1309,
    new_n1310, new_n1311, new_n1312, new_n1313, new_n1314, new_n1315,
    new_n1316, new_n1317, new_n1318, new_n1319, new_n1320, new_n1321,
    new_n1322, new_n1323, new_n1324, new_n1325, new_n1326, new_n1327,
    new_n1328, new_n1329, new_n1330, new_n1331, new_n1332, new_n1333,
    new_n1334, new_n1335, new_n1336, new_n1337, new_n1338, new_n1339,
    new_n1340, new_n1341, new_n1342, new_n1343, new_n1344, new_n1345,
    new_n1346, new_n1347, new_n1348, new_n1349, new_n1351, new_n1352,
    new_n1353, new_n1354, new_n1355, new_n1356, new_n1357, new_n1358,
    new_n1359, new_n1360, new_n1361, new_n1362, new_n1363, new_n1364,
    new_n1365, new_n1366, new_n1367, new_n1368, new_n1369, new_n1370,
    new_n1371, new_n1372, new_n1373, new_n1374, new_n1375, new_n1376,
    new_n1377, new_n1378, new_n1379, new_n1380, new_n1381, new_n1382,
    new_n1383, new_n1384, new_n1385, new_n1386, new_n1387, new_n1388,
    new_n1389, new_n1390, new_n1391, new_n1392, new_n1393, new_n1394,
    new_n1395, new_n1396, new_n1397, new_n1398, new_n1399, new_n1400,
    new_n1401, new_n1402, new_n1403, new_n1404, new_n1405, new_n1406,
    new_n1407, new_n1408, new_n1409, new_n1410, new_n1411, new_n1412,
    new_n1413, new_n1414, new_n1415, new_n1416, new_n1417, new_n1418,
    new_n1419, new_n1420, new_n1421, new_n1422, new_n1423, new_n1424,
    new_n1425, new_n1426, new_n1427, new_n1428, new_n1429, new_n1430,
    new_n1431, new_n1432, new_n1433, new_n1434, new_n1435, new_n1436,
    new_n1437, new_n1438, new_n1439, new_n1440, new_n1441, new_n1442,
    new_n1443, new_n1444, new_n1445, new_n1446, new_n1447, new_n1448,
    new_n1449, new_n1450, new_n1451, new_n1452, new_n1453, new_n1454,
    new_n1455, new_n1456, new_n1457, new_n1458, new_n1459, new_n1460,
    new_n1461, new_n1462, new_n1463, new_n1464, new_n1465, new_n1466,
    new_n1467, new_n1468, new_n1469, new_n1470, new_n1471, new_n1473,
    new_n1474, new_n1475, new_n1476, new_n1477, new_n1478, new_n1479,
    new_n1480, new_n1481, new_n1482, new_n1483, new_n1484, new_n1485,
    new_n1486, new_n1487, new_n1488, new_n1489, new_n1490, new_n1491,
    new_n1492, new_n1493, new_n1494, new_n1495, new_n1496, new_n1497,
    new_n1498, new_n1499, new_n1500, new_n1501, new_n1502, new_n1503,
    new_n1504, new_n1505, new_n1506, new_n1507, new_n1508, new_n1509,
    new_n1510, new_n1511, new_n1512, new_n1513, new_n1514, new_n1515,
    new_n1516, new_n1517, new_n1518, new_n1519, new_n1520, new_n1521,
    new_n1522, new_n1523, new_n1524, new_n1525, new_n1526, new_n1527,
    new_n1528, new_n1529, new_n1530, new_n1531, new_n1532, new_n1533,
    new_n1534, new_n1535, new_n1536, new_n1537, new_n1538, new_n1539,
    new_n1540, new_n1541, new_n1542, new_n1543, new_n1544, new_n1545,
    new_n1546, new_n1547, new_n1548, new_n1549, new_n1550, new_n1551,
    new_n1552, new_n1553, new_n1554, new_n1555, new_n1556, new_n1557,
    new_n1558, new_n1559, new_n1560, new_n1561, new_n1562, new_n1563,
    new_n1564, new_n1565, new_n1566, new_n1567, new_n1568, new_n1569,
    new_n1570, new_n1571, new_n1572, new_n1573, new_n1574, new_n1575,
    new_n1576, new_n1577, new_n1578, new_n1579, new_n1580, new_n1581,
    new_n1582, new_n1583, new_n1584, new_n1585, new_n1586, new_n1587,
    new_n1588, new_n1589, new_n1590, new_n1591, new_n1592, new_n1593,
    new_n1595, new_n1596, new_n1597, new_n1598, new_n1599, new_n1600,
    new_n1601, new_n1602, new_n1603, new_n1604, new_n1605, new_n1606,
    new_n1607, new_n1608, new_n1609, new_n1610, new_n1611, new_n1612,
    new_n1613, new_n1614, new_n1615, new_n1616, new_n1617, new_n1618,
    new_n1619, new_n1620, new_n1621, new_n1622, new_n1623, new_n1624,
    new_n1625, new_n1626, new_n1627, new_n1628, new_n1629, new_n1630,
    new_n1631, new_n1632, new_n1633, new_n1634, new_n1635, new_n1636,
    new_n1637, new_n1638, new_n1639, new_n1640, new_n1641, new_n1642,
    new_n1643, new_n1644, new_n1645, new_n1646, new_n1647, new_n1648,
    new_n1649, new_n1650, new_n1651, new_n1652, new_n1653, new_n1654,
    new_n1655, new_n1656, new_n1657, new_n1658, new_n1659, new_n1660,
    new_n1661, new_n1662, new_n1663, new_n1664, new_n1665, new_n1666,
    new_n1667, new_n1668, new_n1669, new_n1670, new_n1671, new_n1672,
    new_n1673, new_n1674, new_n1675, new_n1676, new_n1677, new_n1678,
    new_n1679, new_n1680, new_n1681, new_n1682, new_n1683, new_n1684,
    new_n1685, new_n1686, new_n1687, new_n1688, new_n1689, new_n1690,
    new_n1691, new_n1692, new_n1693, new_n1694, new_n1695, new_n1696,
    new_n1697, new_n1698, new_n1699, new_n1700, new_n1701, new_n1702,
    new_n1703, new_n1704, new_n1705, new_n1706, new_n1707, new_n1708,
    new_n1709, new_n1710, new_n1711, new_n1712, new_n1713, new_n1714,
    new_n1715, new_n1716, new_n1717, new_n1718, new_n1719, new_n1720,
    new_n1721, new_n1722, new_n1723, new_n1724, new_n1725, new_n1726,
    new_n1727, new_n1728, new_n1729, new_n1730, new_n1732, new_n1733,
    new_n1734, new_n1735, new_n1736, new_n1737, new_n1738, new_n1739,
    new_n1740, new_n1741, new_n1742, new_n1743, new_n1744, new_n1745,
    new_n1746, new_n1747, new_n1748, new_n1749, new_n1750, new_n1751,
    new_n1752, new_n1753, new_n1754, new_n1755, new_n1756, new_n1757,
    new_n1758, new_n1759, new_n1760, new_n1761, new_n1762, new_n1763,
    new_n1764, new_n1765, new_n1766, new_n1767, new_n1768, new_n1769,
    new_n1770, new_n1771, new_n1772, new_n1773, new_n1774, new_n1775,
    new_n1776, new_n1777, new_n1778, new_n1779, new_n1780, new_n1781,
    new_n1782, new_n1783, new_n1784, new_n1785, new_n1786, new_n1787,
    new_n1788, new_n1789, new_n1790, new_n1791, new_n1792, new_n1793,
    new_n1794, new_n1795, new_n1796, new_n1797, new_n1798, new_n1799,
    new_n1800, new_n1801, new_n1802, new_n1803, new_n1804, new_n1805,
    new_n1806, new_n1807, new_n1808, new_n1809, new_n1810, new_n1811,
    new_n1812, new_n1813, new_n1814, new_n1815, new_n1816, new_n1817,
    new_n1818, new_n1819, new_n1820, new_n1821, new_n1822, new_n1823,
    new_n1824, new_n1825, new_n1826, new_n1827, new_n1828, new_n1829,
    new_n1830, new_n1831, new_n1832, new_n1833, new_n1834, new_n1835,
    new_n1836, new_n1837, new_n1838, new_n1839, new_n1840, new_n1841,
    new_n1842, new_n1843, new_n1844, new_n1845, new_n1846, new_n1847,
    new_n1848, new_n1849, new_n1850, new_n1851, new_n1852, new_n1853,
    new_n1854, new_n1855, new_n1856, new_n1857, new_n1858, new_n1859,
    new_n1860, new_n1861, new_n1862, new_n1863, new_n1864, new_n1865,
    new_n1866, new_n1868, new_n1869, new_n1870, new_n1871, new_n1872,
    new_n1873, new_n1874, new_n1875, new_n1876, new_n1877, new_n1878,
    new_n1879, new_n1880, new_n1881, new_n1882, new_n1883, new_n1884,
    new_n1885, new_n1886, new_n1887, new_n1888, new_n1889, new_n1890,
    new_n1891, new_n1892, new_n1893, new_n1894, new_n1895, new_n1896,
    new_n1897, new_n1898, new_n1899, new_n1900, new_n1901, new_n1902,
    new_n1903, new_n1904, new_n1905, new_n1906, new_n1907, new_n1908,
    new_n1909, new_n1910, new_n1911, new_n1912, new_n1913, new_n1914,
    new_n1915, new_n1916, new_n1917, new_n1918, new_n1919, new_n1920,
    new_n1921, new_n1922, new_n1923, new_n1924, new_n1925, new_n1926,
    new_n1927, new_n1928, new_n1929, new_n1930, new_n1931, new_n1932,
    new_n1933, new_n1934, new_n1935, new_n1936, new_n1937, new_n1938,
    new_n1939, new_n1940, new_n1941, new_n1942, new_n1943, new_n1944,
    new_n1945, new_n1946, new_n1947, new_n1948, new_n1949, new_n1950,
    new_n1951, new_n1952, new_n1953, new_n1954, new_n1955, new_n1956,
    new_n1957, new_n1958, new_n1959, new_n1960, new_n1961, new_n1962,
    new_n1963, new_n1964, new_n1965, new_n1966, new_n1967, new_n1968,
    new_n1969, new_n1970, new_n1971, new_n1972, new_n1973, new_n1974,
    new_n1975, new_n1976, new_n1977, new_n1978, new_n1979, new_n1980,
    new_n1981, new_n1982, new_n1983, new_n1984, new_n1985, new_n1986,
    new_n1987, new_n1988, new_n1989, new_n1990, new_n1991, new_n1992,
    new_n1993, new_n1994, new_n1995, new_n1996, new_n1997, new_n1998,
    new_n1999, new_n2000, new_n2001, new_n2002, new_n2003, new_n2004,
    new_n2005, new_n2006, new_n2007, new_n2008, new_n2010, new_n2011,
    new_n2012, new_n2013, new_n2014, new_n2015, new_n2016, new_n2017,
    new_n2018, new_n2019, new_n2020, new_n2021, new_n2022, new_n2023,
    new_n2024, new_n2025, new_n2026, new_n2027, new_n2028, new_n2029,
    new_n2030, new_n2031, new_n2032, new_n2033, new_n2034, new_n2035,
    new_n2036, new_n2037, new_n2038, new_n2039, new_n2040, new_n2041,
    new_n2042, new_n2043, new_n2044, new_n2045, new_n2046, new_n2047,
    new_n2048, new_n2049, new_n2050, new_n2051, new_n2052, new_n2053,
    new_n2054, new_n2055, new_n2056, new_n2057, new_n2058, new_n2059,
    new_n2060, new_n2061, new_n2062, new_n2063, new_n2064, new_n2065,
    new_n2066, new_n2067, new_n2068, new_n2069, new_n2070, new_n2071,
    new_n2072, new_n2073, new_n2074, new_n2075, new_n2076, new_n2077,
    new_n2078, new_n2079, new_n2080, new_n2081, new_n2082, new_n2083,
    new_n2084, new_n2085, new_n2086, new_n2087, new_n2088, new_n2089,
    new_n2090, new_n2091, new_n2092, new_n2093, new_n2094, new_n2095,
    new_n2096, new_n2097, new_n2098, new_n2099, new_n2100, new_n2101,
    new_n2102, new_n2103, new_n2104, new_n2105, new_n2106, new_n2107,
    new_n2108, new_n2109, new_n2110, new_n2111, new_n2112, new_n2113,
    new_n2114, new_n2115, new_n2116, new_n2117, new_n2118, new_n2119,
    new_n2120, new_n2121, new_n2122, new_n2123, new_n2124, new_n2125,
    new_n2126, new_n2127, new_n2128, new_n2129, new_n2130, new_n2131,
    new_n2132, new_n2133, new_n2134, new_n2135, new_n2136, new_n2137,
    new_n2138, new_n2139, new_n2140, new_n2141, new_n2142, new_n2143,
    new_n2144, new_n2145, new_n2146, new_n2147, new_n2148, new_n2149,
    new_n2150, new_n2151, new_n2152, new_n2153, new_n2154, new_n2155,
    new_n2156, new_n2157, new_n2158, new_n2159, new_n2161, new_n2162,
    new_n2163, new_n2164, new_n2165, new_n2166, new_n2167, new_n2168,
    new_n2169, new_n2170, new_n2171, new_n2172, new_n2173, new_n2174,
    new_n2175, new_n2176, new_n2177, new_n2178, new_n2179, new_n2180,
    new_n2181, new_n2182, new_n2183, new_n2184, new_n2185, new_n2186,
    new_n2187, new_n2188, new_n2189, new_n2190, new_n2191, new_n2192,
    new_n2193, new_n2194, new_n2195, new_n2196, new_n2197, new_n2198,
    new_n2199, new_n2200, new_n2201, new_n2202, new_n2203, new_n2204,
    new_n2205, new_n2206, new_n2207, new_n2208, new_n2209, new_n2210,
    new_n2211, new_n2212, new_n2213, new_n2214, new_n2215, new_n2216,
    new_n2217, new_n2218, new_n2219, new_n2220, new_n2221, new_n2222,
    new_n2223, new_n2224, new_n2225, new_n2226, new_n2227, new_n2228,
    new_n2229, new_n2230, new_n2231, new_n2232, new_n2233, new_n2234,
    new_n2235, new_n2236, new_n2237, new_n2238, new_n2239, new_n2240,
    new_n2241, new_n2242, new_n2243, new_n2244, new_n2245, new_n2246,
    new_n2247, new_n2248, new_n2249, new_n2250, new_n2251, new_n2252,
    new_n2253, new_n2254, new_n2255, new_n2256, new_n2257, new_n2258,
    new_n2259, new_n2260, new_n2261, new_n2262, new_n2263, new_n2264,
    new_n2265, new_n2266, new_n2267, new_n2268, new_n2269, new_n2270,
    new_n2271, new_n2272, new_n2273, new_n2274, new_n2275, new_n2276,
    new_n2277, new_n2278, new_n2279, new_n2280, new_n2281, new_n2282,
    new_n2283, new_n2284, new_n2285, new_n2286, new_n2287, new_n2288,
    new_n2289, new_n2290, new_n2291, new_n2292, new_n2293, new_n2294,
    new_n2295, new_n2296, new_n2297, new_n2298, new_n2299, new_n2300,
    new_n2301, new_n2302, new_n2303, new_n2304, new_n2305, new_n2306,
    new_n2307, new_n2308, new_n2309, new_n2310, new_n2311, new_n2312,
    new_n2313, new_n2314, new_n2315, new_n2316, new_n2317, new_n2319,
    new_n2320, new_n2321, new_n2322, new_n2323, new_n2324, new_n2325,
    new_n2326, new_n2327, new_n2328, new_n2329, new_n2330, new_n2331,
    new_n2332, new_n2333, new_n2334, new_n2335, new_n2336, new_n2337,
    new_n2338, new_n2339, new_n2340, new_n2341, new_n2342, new_n2343,
    new_n2344, new_n2345, new_n2346, new_n2347, new_n2348, new_n2349,
    new_n2350, new_n2351, new_n2352, new_n2353, new_n2354, new_n2355,
    new_n2356, new_n2357, new_n2358, new_n2359, new_n2360, new_n2361,
    new_n2362, new_n2363, new_n2364, new_n2365, new_n2366, new_n2367,
    new_n2368, new_n2369, new_n2370, new_n2371, new_n2372, new_n2373,
    new_n2374, new_n2375, new_n2376, new_n2377, new_n2378, new_n2379,
    new_n2380, new_n2381, new_n2382, new_n2383, new_n2384, new_n2385,
    new_n2386, new_n2387, new_n2388, new_n2389, new_n2390, new_n2391,
    new_n2392, new_n2393, new_n2394, new_n2395, new_n2396, new_n2397,
    new_n2398, new_n2399, new_n2400, new_n2401, new_n2402, new_n2403,
    new_n2404, new_n2405, new_n2406, new_n2407, new_n2408, new_n2409,
    new_n2410, new_n2411, new_n2412, new_n2413, new_n2414, new_n2415,
    new_n2416, new_n2417, new_n2418, new_n2419, new_n2420, new_n2421,
    new_n2422, new_n2423, new_n2424, new_n2425, new_n2426, new_n2427,
    new_n2428, new_n2429, new_n2430, new_n2431, new_n2432, new_n2433,
    new_n2434, new_n2435, new_n2436, new_n2437, new_n2438, new_n2439,
    new_n2440, new_n2441, new_n2442, new_n2443, new_n2444, new_n2445,
    new_n2446, new_n2447, new_n2448, new_n2449, new_n2450, new_n2451,
    new_n2452, new_n2453, new_n2454, new_n2455, new_n2456, new_n2457,
    new_n2458, new_n2459, new_n2460, new_n2461, new_n2462, new_n2463,
    new_n2464, new_n2465, new_n2466, new_n2467, new_n2468, new_n2469,
    new_n2470, new_n2471, new_n2472, new_n2473, new_n2474, new_n2475,
    new_n2476, new_n2477, new_n2478, new_n2480, new_n2481, new_n2482,
    new_n2483, new_n2484, new_n2485, new_n2486, new_n2487, new_n2488,
    new_n2489, new_n2490, new_n2491, new_n2492, new_n2493, new_n2494,
    new_n2495, new_n2496, new_n2497, new_n2498, new_n2499, new_n2500,
    new_n2501, new_n2502, new_n2503, new_n2504, new_n2505, new_n2506,
    new_n2507, new_n2508, new_n2509, new_n2510, new_n2511, new_n2512,
    new_n2513, new_n2514, new_n2515, new_n2516, new_n2517, new_n2518,
    new_n2519, new_n2520, new_n2521, new_n2522, new_n2523, new_n2524,
    new_n2525, new_n2526, new_n2527, new_n2528, new_n2529, new_n2530,
    new_n2531, new_n2532, new_n2533, new_n2534, new_n2535, new_n2536,
    new_n2537, new_n2538, new_n2539, new_n2540, new_n2541, new_n2542,
    new_n2543, new_n2544, new_n2545, new_n2546, new_n2547, new_n2548,
    new_n2549, new_n2550, new_n2551, new_n2552, new_n2553, new_n2554,
    new_n2555, new_n2556, new_n2557, new_n2558, new_n2559, new_n2560,
    new_n2561, new_n2562, new_n2563, new_n2564, new_n2565, new_n2566,
    new_n2567, new_n2568, new_n2569, new_n2570, new_n2571, new_n2572,
    new_n2573, new_n2574, new_n2575, new_n2576, new_n2577, new_n2578,
    new_n2579, new_n2580, new_n2581, new_n2582, new_n2583, new_n2584,
    new_n2585, new_n2586, new_n2587, new_n2588, new_n2589, new_n2590,
    new_n2591, new_n2592, new_n2593, new_n2594, new_n2595, new_n2596,
    new_n2597, new_n2598, new_n2599, new_n2600, new_n2601, new_n2602,
    new_n2603, new_n2604, new_n2605, new_n2606, new_n2607, new_n2608,
    new_n2609, new_n2610, new_n2611, new_n2612, new_n2613, new_n2614,
    new_n2615, new_n2616, new_n2617, new_n2618, new_n2619, new_n2620,
    new_n2621, new_n2622, new_n2623, new_n2624, new_n2625, new_n2626,
    new_n2627, new_n2628, new_n2629, new_n2630, new_n2631, new_n2632,
    new_n2633, new_n2634, new_n2635, new_n2636, new_n2637, new_n2638,
    new_n2639, new_n2640, new_n2641, new_n2642, new_n2643, new_n2644,
    new_n2645, new_n2646, new_n2648, new_n2649, new_n2650, new_n2651,
    new_n2652, new_n2653, new_n2654, new_n2655, new_n2656, new_n2657,
    new_n2658, new_n2659, new_n2660, new_n2661, new_n2662, new_n2663,
    new_n2664, new_n2665, new_n2666, new_n2667, new_n2668, new_n2669,
    new_n2670, new_n2671, new_n2672, new_n2673, new_n2674, new_n2675,
    new_n2676, new_n2677, new_n2678, new_n2679, new_n2680, new_n2681,
    new_n2682, new_n2683, new_n2684, new_n2685, new_n2686, new_n2687,
    new_n2688, new_n2689, new_n2690, new_n2691, new_n2692, new_n2693,
    new_n2694, new_n2695, new_n2696, new_n2697, new_n2698, new_n2699,
    new_n2700, new_n2701, new_n2702, new_n2703, new_n2704, new_n2705,
    new_n2706, new_n2707, new_n2708, new_n2709, new_n2710, new_n2711,
    new_n2712, new_n2713, new_n2714, new_n2715, new_n2716, new_n2717,
    new_n2718, new_n2719, new_n2720, new_n2721, new_n2722, new_n2723,
    new_n2724, new_n2725, new_n2726, new_n2727, new_n2728, new_n2729,
    new_n2730, new_n2731, new_n2732, new_n2733, new_n2734, new_n2735,
    new_n2736, new_n2737, new_n2738, new_n2739, new_n2740, new_n2741,
    new_n2742, new_n2743, new_n2744, new_n2745, new_n2746, new_n2747,
    new_n2748, new_n2749, new_n2750, new_n2751, new_n2752, new_n2753,
    new_n2754, new_n2755, new_n2756, new_n2757, new_n2758, new_n2759,
    new_n2760, new_n2761, new_n2762, new_n2763, new_n2764, new_n2765,
    new_n2766, new_n2767, new_n2768, new_n2769, new_n2770, new_n2771,
    new_n2772, new_n2773, new_n2774, new_n2775, new_n2776, new_n2777,
    new_n2778, new_n2779, new_n2780, new_n2781, new_n2782, new_n2783,
    new_n2784, new_n2785, new_n2786, new_n2787, new_n2788, new_n2789,
    new_n2790, new_n2791, new_n2792, new_n2793, new_n2794, new_n2795,
    new_n2796, new_n2797, new_n2798, new_n2799, new_n2800, new_n2801,
    new_n2802, new_n2803, new_n2804, new_n2805, new_n2806, new_n2807,
    new_n2808, new_n2809, new_n2810, new_n2811, new_n2812, new_n2813,
    new_n2814, new_n2815, new_n2816, new_n2817, new_n2818, new_n2819,
    new_n2820, new_n2822, new_n2823, new_n2824, new_n2825, new_n2826,
    new_n2827, new_n2828, new_n2829, new_n2830, new_n2831, new_n2832,
    new_n2833, new_n2834, new_n2835, new_n2836, new_n2837, new_n2838,
    new_n2839, new_n2840, new_n2841, new_n2842, new_n2843, new_n2844,
    new_n2845, new_n2846, new_n2847, new_n2848, new_n2849, new_n2850,
    new_n2851, new_n2852, new_n2853, new_n2854, new_n2855, new_n2856,
    new_n2857, new_n2858, new_n2859, new_n2860, new_n2861, new_n2862,
    new_n2863, new_n2864, new_n2865, new_n2866, new_n2867, new_n2868,
    new_n2869, new_n2870, new_n2871, new_n2872, new_n2873, new_n2874,
    new_n2875, new_n2876, new_n2877, new_n2878, new_n2879, new_n2880,
    new_n2881, new_n2882, new_n2883, new_n2884, new_n2885, new_n2886,
    new_n2887, new_n2888, new_n2889, new_n2890, new_n2891, new_n2892,
    new_n2893, new_n2894, new_n2895, new_n2896, new_n2897, new_n2898,
    new_n2899, new_n2900, new_n2901, new_n2902, new_n2903, new_n2904,
    new_n2905, new_n2906, new_n2907, new_n2908, new_n2909, new_n2910,
    new_n2911, new_n2912, new_n2913, new_n2914, new_n2915, new_n2916,
    new_n2917, new_n2918, new_n2919, new_n2920, new_n2921, new_n2922,
    new_n2923, new_n2924, new_n2925, new_n2926, new_n2927, new_n2928,
    new_n2929, new_n2930, new_n2931, new_n2932, new_n2933, new_n2934,
    new_n2935, new_n2936, new_n2937, new_n2938, new_n2939, new_n2940,
    new_n2941, new_n2942, new_n2943, new_n2944, new_n2945, new_n2946,
    new_n2947, new_n2948, new_n2949, new_n2950, new_n2951, new_n2952,
    new_n2953, new_n2954, new_n2955, new_n2956, new_n2957, new_n2958,
    new_n2959, new_n2960, new_n2961, new_n2962, new_n2963, new_n2964,
    new_n2965, new_n2966, new_n2967, new_n2968, new_n2969, new_n2970,
    new_n2971, new_n2972, new_n2973, new_n2974, new_n2975, new_n2976,
    new_n2977, new_n2978, new_n2979, new_n2980, new_n2981, new_n2982,
    new_n2983, new_n2984, new_n2985, new_n2986, new_n2987, new_n2988,
    new_n2989, new_n2990, new_n2991, new_n2992, new_n2993, new_n2994,
    new_n2995, new_n2996, new_n2997, new_n2998, new_n2999, new_n3000,
    new_n3001, new_n3003, new_n3004, new_n3005, new_n3006, new_n3007,
    new_n3008, new_n3009, new_n3010, new_n3011, new_n3012, new_n3013,
    new_n3014, new_n3015, new_n3016, new_n3017, new_n3018, new_n3019,
    new_n3020, new_n3021, new_n3022, new_n3023, new_n3024, new_n3025,
    new_n3026, new_n3027, new_n3028, new_n3029, new_n3030, new_n3031,
    new_n3032, new_n3033, new_n3034, new_n3035, new_n3036, new_n3037,
    new_n3038, new_n3039, new_n3040, new_n3041, new_n3042, new_n3043,
    new_n3044, new_n3045, new_n3046, new_n3047, new_n3048, new_n3049,
    new_n3050, new_n3051, new_n3052, new_n3053, new_n3054, new_n3055,
    new_n3056, new_n3057, new_n3058, new_n3059, new_n3060, new_n3061,
    new_n3062, new_n3063, new_n3064, new_n3065, new_n3066, new_n3067,
    new_n3068, new_n3069, new_n3070, new_n3071, new_n3072, new_n3073,
    new_n3074, new_n3075, new_n3076, new_n3077, new_n3078, new_n3079,
    new_n3080, new_n3081, new_n3082, new_n3083, new_n3084, new_n3085,
    new_n3086, new_n3087, new_n3088, new_n3089, new_n3090, new_n3091,
    new_n3092, new_n3093, new_n3094, new_n3095, new_n3096, new_n3097,
    new_n3098, new_n3099, new_n3100, new_n3101, new_n3102, new_n3103,
    new_n3104, new_n3105, new_n3106, new_n3107, new_n3108, new_n3109,
    new_n3110, new_n3111, new_n3112, new_n3113, new_n3114, new_n3115,
    new_n3116, new_n3117, new_n3118, new_n3119, new_n3120, new_n3121,
    new_n3122, new_n3123, new_n3124, new_n3125, new_n3126, new_n3127,
    new_n3128, new_n3129, new_n3130, new_n3131, new_n3132, new_n3133,
    new_n3134, new_n3135, new_n3136, new_n3137, new_n3138, new_n3139,
    new_n3140, new_n3141, new_n3142, new_n3143, new_n3144, new_n3145,
    new_n3146, new_n3147, new_n3148, new_n3149, new_n3150, new_n3151,
    new_n3152, new_n3153, new_n3154, new_n3155, new_n3156, new_n3157,
    new_n3158, new_n3159, new_n3160, new_n3161, new_n3162, new_n3163,
    new_n3164, new_n3165, new_n3166, new_n3167, new_n3168, new_n3169,
    new_n3170, new_n3171, new_n3172, new_n3173, new_n3174, new_n3175,
    new_n3176, new_n3177, new_n3178, new_n3179, new_n3180, new_n3181,
    new_n3182, new_n3183, new_n3184, new_n3185, new_n3186, new_n3188,
    new_n3189, new_n3190, new_n3191, new_n3192, new_n3193, new_n3194,
    new_n3195, new_n3196, new_n3197, new_n3198, new_n3199, new_n3200,
    new_n3201, new_n3202, new_n3203, new_n3204, new_n3205, new_n3206,
    new_n3207, new_n3208, new_n3209, new_n3210, new_n3211, new_n3212,
    new_n3213, new_n3214, new_n3215, new_n3216, new_n3217, new_n3218,
    new_n3219, new_n3220, new_n3221, new_n3222, new_n3223, new_n3224,
    new_n3225, new_n3226, new_n3227, new_n3228, new_n3229, new_n3230,
    new_n3231, new_n3232, new_n3233, new_n3234, new_n3235, new_n3236,
    new_n3237, new_n3238, new_n3239, new_n3240, new_n3241, new_n3242,
    new_n3243, new_n3244, new_n3245, new_n3246, new_n3247, new_n3248,
    new_n3249, new_n3250, new_n3251, new_n3252, new_n3253, new_n3254,
    new_n3255, new_n3256, new_n3257, new_n3258, new_n3259, new_n3260,
    new_n3261, new_n3262, new_n3263, new_n3264, new_n3265, new_n3266,
    new_n3267, new_n3268, new_n3269, new_n3270, new_n3271, new_n3272,
    new_n3273, new_n3274, new_n3275, new_n3276, new_n3277, new_n3278,
    new_n3279, new_n3280, new_n3281, new_n3282, new_n3283, new_n3284,
    new_n3285, new_n3286, new_n3287, new_n3288, new_n3289, new_n3290,
    new_n3291, new_n3292, new_n3293, new_n3294, new_n3295, new_n3296,
    new_n3297, new_n3298, new_n3299, new_n3300, new_n3301, new_n3302,
    new_n3303, new_n3304, new_n3305, new_n3306, new_n3307, new_n3308,
    new_n3309, new_n3310, new_n3311, new_n3312, new_n3313, new_n3314,
    new_n3315, new_n3316, new_n3317, new_n3318, new_n3319, new_n3320,
    new_n3321, new_n3322, new_n3323, new_n3324, new_n3325, new_n3326,
    new_n3327, new_n3328, new_n3329, new_n3330, new_n3331, new_n3332,
    new_n3333, new_n3334, new_n3335, new_n3336, new_n3337, new_n3338,
    new_n3339, new_n3340, new_n3341, new_n3342, new_n3343, new_n3344,
    new_n3345, new_n3346, new_n3347, new_n3348, new_n3349, new_n3350,
    new_n3351, new_n3352, new_n3353, new_n3354, new_n3355, new_n3356,
    new_n3357, new_n3358, new_n3359, new_n3360, new_n3361, new_n3362,
    new_n3363, new_n3364, new_n3365, new_n3366, new_n3367, new_n3368,
    new_n3369, new_n3370, new_n3371, new_n3372, new_n3373, new_n3374,
    new_n3375, new_n3376, new_n3377, new_n3378, new_n3379, new_n3381,
    new_n3382, new_n3383, new_n3384, new_n3385, new_n3386, new_n3387,
    new_n3388, new_n3389, new_n3390, new_n3391, new_n3392, new_n3393,
    new_n3394, new_n3395, new_n3396, new_n3397, new_n3398, new_n3399,
    new_n3400, new_n3401, new_n3402, new_n3403, new_n3404, new_n3405,
    new_n3406, new_n3407, new_n3408, new_n3409, new_n3410, new_n3411,
    new_n3412, new_n3413, new_n3414, new_n3415, new_n3416, new_n3417,
    new_n3418, new_n3419, new_n3420, new_n3421, new_n3422, new_n3423,
    new_n3424, new_n3425, new_n3426, new_n3427, new_n3428, new_n3429,
    new_n3430, new_n3431, new_n3432, new_n3433, new_n3434, new_n3435,
    new_n3436, new_n3437, new_n3438, new_n3439, new_n3440, new_n3441,
    new_n3442, new_n3443, new_n3444, new_n3445, new_n3446, new_n3447,
    new_n3448, new_n3449, new_n3450, new_n3451, new_n3452, new_n3453,
    new_n3454, new_n3455, new_n3456, new_n3457, new_n3458, new_n3459,
    new_n3460, new_n3461, new_n3462, new_n3463, new_n3464, new_n3465,
    new_n3466, new_n3467, new_n3468, new_n3469, new_n3470, new_n3471,
    new_n3472, new_n3473, new_n3474, new_n3475, new_n3476, new_n3477,
    new_n3478, new_n3479, new_n3480, new_n3481, new_n3482, new_n3483,
    new_n3484, new_n3485, new_n3486, new_n3487, new_n3488, new_n3489,
    new_n3490, new_n3491, new_n3492, new_n3493, new_n3494, new_n3495,
    new_n3496, new_n3497, new_n3498, new_n3499, new_n3500, new_n3501,
    new_n3502, new_n3503, new_n3504, new_n3505, new_n3506, new_n3507,
    new_n3508, new_n3509, new_n3510, new_n3511, new_n3512, new_n3513,
    new_n3514, new_n3515, new_n3516, new_n3517, new_n3518, new_n3519,
    new_n3520, new_n3521, new_n3522, new_n3523, new_n3524, new_n3525,
    new_n3526, new_n3527, new_n3528, new_n3529, new_n3530, new_n3531,
    new_n3532, new_n3533, new_n3534, new_n3535, new_n3536, new_n3537,
    new_n3538, new_n3539, new_n3540, new_n3541, new_n3542, new_n3543,
    new_n3544, new_n3545, new_n3546, new_n3547, new_n3548, new_n3549,
    new_n3550, new_n3551, new_n3552, new_n3553, new_n3554, new_n3555,
    new_n3556, new_n3557, new_n3558, new_n3559, new_n3560, new_n3561,
    new_n3562, new_n3563, new_n3564, new_n3565, new_n3566, new_n3567,
    new_n3568, new_n3569, new_n3570, new_n3571, new_n3572, new_n3573,
    new_n3575, new_n3576, new_n3577, new_n3578, new_n3579, new_n3580,
    new_n3581, new_n3582, new_n3583, new_n3584, new_n3585, new_n3586,
    new_n3587, new_n3588, new_n3589, new_n3590, new_n3591, new_n3592,
    new_n3593, new_n3594, new_n3595, new_n3596, new_n3597, new_n3598,
    new_n3599, new_n3600, new_n3601, new_n3602, new_n3603, new_n3604,
    new_n3605, new_n3606, new_n3607, new_n3608, new_n3609, new_n3610,
    new_n3611, new_n3612, new_n3613, new_n3614, new_n3615, new_n3616,
    new_n3617, new_n3618, new_n3619, new_n3620, new_n3621, new_n3622,
    new_n3623, new_n3624, new_n3625, new_n3626, new_n3627, new_n3628,
    new_n3629, new_n3630, new_n3631, new_n3632, new_n3633, new_n3634,
    new_n3635, new_n3636, new_n3637, new_n3638, new_n3639, new_n3640,
    new_n3641, new_n3642, new_n3643, new_n3644, new_n3645, new_n3646,
    new_n3647, new_n3648, new_n3649, new_n3650, new_n3651, new_n3652,
    new_n3653, new_n3654, new_n3655, new_n3656, new_n3657, new_n3658,
    new_n3659, new_n3660, new_n3661, new_n3662, new_n3663, new_n3664,
    new_n3665, new_n3666, new_n3667, new_n3668, new_n3669, new_n3670,
    new_n3671, new_n3672, new_n3673, new_n3674, new_n3675, new_n3676,
    new_n3677, new_n3678, new_n3679, new_n3680, new_n3681, new_n3682,
    new_n3683, new_n3684, new_n3685, new_n3686, new_n3687, new_n3688,
    new_n3689, new_n3690, new_n3691, new_n3692, new_n3693, new_n3694,
    new_n3695, new_n3696, new_n3697, new_n3698, new_n3699, new_n3700,
    new_n3701, new_n3702, new_n3703, new_n3704, new_n3705, new_n3706,
    new_n3707, new_n3708, new_n3709, new_n3710, new_n3711, new_n3712,
    new_n3713, new_n3714, new_n3715, new_n3716, new_n3717, new_n3718,
    new_n3719, new_n3720, new_n3721, new_n3722, new_n3723, new_n3724,
    new_n3725, new_n3726, new_n3727, new_n3728, new_n3729, new_n3730,
    new_n3731, new_n3732, new_n3733, new_n3734, new_n3735, new_n3736,
    new_n3737, new_n3738, new_n3739, new_n3740, new_n3741, new_n3742,
    new_n3743, new_n3744, new_n3745, new_n3746, new_n3747, new_n3748,
    new_n3749, new_n3750, new_n3751, new_n3752, new_n3753, new_n3754,
    new_n3755, new_n3756, new_n3757, new_n3758, new_n3759, new_n3760,
    new_n3761, new_n3762, new_n3763, new_n3764, new_n3765, new_n3766,
    new_n3767, new_n3768, new_n3769, new_n3770, new_n3771, new_n3772,
    new_n3773, new_n3774, new_n3775, new_n3776, new_n3777, new_n3778,
    new_n3779, new_n3780, new_n3782, new_n3783, new_n3784, new_n3785,
    new_n3786, new_n3787, new_n3788, new_n3789, new_n3790, new_n3791,
    new_n3792, new_n3793, new_n3794, new_n3795, new_n3796, new_n3797,
    new_n3798, new_n3799, new_n3800, new_n3801, new_n3802, new_n3803,
    new_n3804, new_n3805, new_n3806, new_n3807, new_n3808, new_n3809,
    new_n3810, new_n3811, new_n3812, new_n3813, new_n3814, new_n3815,
    new_n3816, new_n3817, new_n3818, new_n3819, new_n3820, new_n3821,
    new_n3822, new_n3823, new_n3824, new_n3825, new_n3826, new_n3827,
    new_n3828, new_n3829, new_n3830, new_n3831, new_n3832, new_n3833,
    new_n3834, new_n3835, new_n3836, new_n3837, new_n3838, new_n3839,
    new_n3840, new_n3841, new_n3842, new_n3843, new_n3844, new_n3845,
    new_n3846, new_n3847, new_n3848, new_n3849, new_n3850, new_n3851,
    new_n3852, new_n3853, new_n3854, new_n3855, new_n3856, new_n3857,
    new_n3858, new_n3859, new_n3860, new_n3861, new_n3862, new_n3863,
    new_n3864, new_n3865, new_n3866, new_n3867, new_n3868, new_n3869,
    new_n3870, new_n3871, new_n3872, new_n3873, new_n3874, new_n3875,
    new_n3876, new_n3877, new_n3878, new_n3879, new_n3880, new_n3881,
    new_n3882, new_n3883, new_n3884, new_n3885, new_n3886, new_n3887,
    new_n3888, new_n3889, new_n3890, new_n3891, new_n3892, new_n3893,
    new_n3894, new_n3895, new_n3896, new_n3897, new_n3898, new_n3899,
    new_n3900, new_n3901, new_n3902, new_n3903, new_n3904, new_n3905,
    new_n3906, new_n3907, new_n3908, new_n3909, new_n3910, new_n3911,
    new_n3912, new_n3913, new_n3914, new_n3915, new_n3916, new_n3917,
    new_n3918, new_n3919, new_n3920, new_n3921, new_n3922, new_n3923,
    new_n3924, new_n3925, new_n3926, new_n3927, new_n3928, new_n3929,
    new_n3930, new_n3931, new_n3932, new_n3933, new_n3934, new_n3935,
    new_n3936, new_n3937, new_n3938, new_n3939, new_n3940, new_n3941,
    new_n3942, new_n3943, new_n3944, new_n3945, new_n3946, new_n3947,
    new_n3948, new_n3949, new_n3950, new_n3951, new_n3952, new_n3953,
    new_n3954, new_n3955, new_n3956, new_n3957, new_n3958, new_n3959,
    new_n3960, new_n3961, new_n3962, new_n3963, new_n3964, new_n3965,
    new_n3966, new_n3967, new_n3968, new_n3969, new_n3970, new_n3971,
    new_n3972, new_n3973, new_n3974, new_n3975, new_n3976, new_n3977,
    new_n3978, new_n3979, new_n3980, new_n3981, new_n3982, new_n3983,
    new_n3984, new_n3985, new_n3987, new_n3988, new_n3989, new_n3990,
    new_n3991, new_n3992, new_n3993, new_n3994, new_n3995, new_n3996,
    new_n3997, new_n3998, new_n3999, new_n4000, new_n4001, new_n4002,
    new_n4003, new_n4004, new_n4005, new_n4006, new_n4007, new_n4008,
    new_n4009, new_n4010, new_n4011, new_n4012, new_n4013, new_n4014,
    new_n4015, new_n4016, new_n4017, new_n4018, new_n4019, new_n4020,
    new_n4021, new_n4022, new_n4023, new_n4024, new_n4025, new_n4026,
    new_n4027, new_n4028, new_n4029, new_n4030, new_n4031, new_n4032,
    new_n4033, new_n4034, new_n4035, new_n4036, new_n4037, new_n4038,
    new_n4039, new_n4040, new_n4041, new_n4042, new_n4043, new_n4044,
    new_n4045, new_n4046, new_n4047, new_n4048, new_n4049, new_n4050,
    new_n4051, new_n4052, new_n4053, new_n4054, new_n4055, new_n4056,
    new_n4057, new_n4058, new_n4059, new_n4060, new_n4061, new_n4062,
    new_n4063, new_n4064, new_n4065, new_n4066, new_n4067, new_n4068,
    new_n4069, new_n4070, new_n4071, new_n4072, new_n4073, new_n4074,
    new_n4075, new_n4076, new_n4077, new_n4078, new_n4079, new_n4080,
    new_n4081, new_n4082, new_n4083, new_n4084, new_n4085, new_n4086,
    new_n4087, new_n4088, new_n4089, new_n4090, new_n4091, new_n4092,
    new_n4093, new_n4094, new_n4095, new_n4096, new_n4097, new_n4098,
    new_n4099, new_n4100, new_n4101, new_n4102, new_n4103, new_n4104,
    new_n4105, new_n4106, new_n4107, new_n4108, new_n4109, new_n4110,
    new_n4111, new_n4112, new_n4113, new_n4114, new_n4115, new_n4116,
    new_n4117, new_n4118, new_n4119, new_n4120, new_n4121, new_n4122,
    new_n4123, new_n4124, new_n4125, new_n4126, new_n4127, new_n4128,
    new_n4129, new_n4130, new_n4131, new_n4132, new_n4133, new_n4134,
    new_n4135, new_n4136, new_n4137, new_n4138, new_n4139, new_n4140,
    new_n4141, new_n4142, new_n4143, new_n4144, new_n4145, new_n4146,
    new_n4147, new_n4148, new_n4149, new_n4150, new_n4151, new_n4152,
    new_n4153, new_n4154, new_n4155, new_n4156, new_n4157, new_n4158,
    new_n4159, new_n4160, new_n4161, new_n4162, new_n4163, new_n4164,
    new_n4165, new_n4166, new_n4167, new_n4168, new_n4169, new_n4170,
    new_n4171, new_n4172, new_n4173, new_n4174, new_n4175, new_n4176,
    new_n4177, new_n4178, new_n4179, new_n4180, new_n4181, new_n4182,
    new_n4183, new_n4184, new_n4185, new_n4186, new_n4187, new_n4188,
    new_n4189, new_n4190, new_n4191, new_n4192, new_n4193, new_n4194,
    new_n4195, new_n4196, new_n4197, new_n4198, new_n4200, new_n4201,
    new_n4202, new_n4203, new_n4204, new_n4205, new_n4206, new_n4207,
    new_n4208, new_n4209, new_n4210, new_n4211, new_n4212, new_n4213,
    new_n4214, new_n4215, new_n4216, new_n4217, new_n4218, new_n4219,
    new_n4220, new_n4221, new_n4222, new_n4223, new_n4224, new_n4225,
    new_n4226, new_n4227, new_n4228, new_n4229, new_n4230, new_n4231,
    new_n4232, new_n4233, new_n4234, new_n4235, new_n4236, new_n4237,
    new_n4238, new_n4239, new_n4240, new_n4241, new_n4242, new_n4243,
    new_n4244, new_n4245, new_n4246, new_n4247, new_n4248, new_n4249,
    new_n4250, new_n4251, new_n4252, new_n4253, new_n4254, new_n4255,
    new_n4256, new_n4257, new_n4258, new_n4259, new_n4260, new_n4261,
    new_n4262, new_n4263, new_n4264, new_n4265, new_n4266, new_n4267,
    new_n4268, new_n4269, new_n4270, new_n4271, new_n4272, new_n4273,
    new_n4274, new_n4275, new_n4276, new_n4277, new_n4278, new_n4279,
    new_n4280, new_n4281, new_n4282, new_n4283, new_n4284, new_n4285,
    new_n4286, new_n4287, new_n4288, new_n4289, new_n4290, new_n4291,
    new_n4292, new_n4293, new_n4294, new_n4295, new_n4296, new_n4297,
    new_n4298, new_n4299, new_n4300, new_n4301, new_n4302, new_n4303,
    new_n4304, new_n4305, new_n4306, new_n4307, new_n4308, new_n4309,
    new_n4310, new_n4311, new_n4312, new_n4313, new_n4314, new_n4315,
    new_n4316, new_n4317, new_n4318, new_n4319, new_n4320, new_n4321,
    new_n4322, new_n4323, new_n4324, new_n4325, new_n4326, new_n4327,
    new_n4328, new_n4329, new_n4330, new_n4331, new_n4332, new_n4333,
    new_n4334, new_n4335, new_n4336, new_n4337, new_n4338, new_n4339,
    new_n4340, new_n4341, new_n4342, new_n4343, new_n4344, new_n4345,
    new_n4346, new_n4347, new_n4348, new_n4349, new_n4350, new_n4351,
    new_n4352, new_n4353, new_n4354, new_n4355, new_n4356, new_n4357,
    new_n4358, new_n4359, new_n4360, new_n4361, new_n4362, new_n4363,
    new_n4364, new_n4365, new_n4366, new_n4367, new_n4368, new_n4369,
    new_n4370, new_n4371, new_n4372, new_n4373, new_n4374, new_n4375,
    new_n4376, new_n4377, new_n4378, new_n4379, new_n4380, new_n4381,
    new_n4382, new_n4383, new_n4384, new_n4385, new_n4386, new_n4387,
    new_n4388, new_n4389, new_n4390, new_n4391, new_n4392, new_n4393,
    new_n4394, new_n4395, new_n4396, new_n4397, new_n4398, new_n4399,
    new_n4400, new_n4401, new_n4402, new_n4403, new_n4404, new_n4405,
    new_n4406, new_n4407, new_n4408, new_n4409, new_n4410, new_n4411,
    new_n4412, new_n4413, new_n4414, new_n4415, new_n4416, new_n4418,
    new_n4419, new_n4420, new_n4421, new_n4422, new_n4423, new_n4424,
    new_n4425, new_n4426, new_n4427, new_n4428, new_n4429, new_n4430,
    new_n4431, new_n4432, new_n4433, new_n4434, new_n4435, new_n4436,
    new_n4437, new_n4438, new_n4439, new_n4440, new_n4441, new_n4442,
    new_n4443, new_n4444, new_n4445, new_n4446, new_n4447, new_n4448,
    new_n4449, new_n4450, new_n4451, new_n4452, new_n4453, new_n4454,
    new_n4455, new_n4456, new_n4457, new_n4458, new_n4459, new_n4460,
    new_n4461, new_n4462, new_n4463, new_n4464, new_n4465, new_n4466,
    new_n4467, new_n4468, new_n4469, new_n4470, new_n4471, new_n4472,
    new_n4473, new_n4474, new_n4475, new_n4476, new_n4477, new_n4478,
    new_n4479, new_n4480, new_n4481, new_n4482, new_n4483, new_n4484,
    new_n4485, new_n4486, new_n4487, new_n4488, new_n4489, new_n4490,
    new_n4491, new_n4492, new_n4493, new_n4494, new_n4495, new_n4496,
    new_n4497, new_n4498, new_n4499, new_n4500, new_n4501, new_n4502,
    new_n4503, new_n4504, new_n4505, new_n4506, new_n4507, new_n4508,
    new_n4509, new_n4510, new_n4511, new_n4512, new_n4513, new_n4514,
    new_n4515, new_n4516, new_n4517, new_n4518, new_n4519, new_n4520,
    new_n4521, new_n4522, new_n4523, new_n4524, new_n4525, new_n4526,
    new_n4527, new_n4528, new_n4529, new_n4530, new_n4531, new_n4532,
    new_n4533, new_n4534, new_n4535, new_n4536, new_n4537, new_n4538,
    new_n4539, new_n4540, new_n4541, new_n4542, new_n4543, new_n4544,
    new_n4545, new_n4546, new_n4547, new_n4548, new_n4549, new_n4550,
    new_n4551, new_n4552, new_n4553, new_n4554, new_n4555, new_n4556,
    new_n4557, new_n4558, new_n4559, new_n4560, new_n4561, new_n4562,
    new_n4563, new_n4564, new_n4565, new_n4566, new_n4567, new_n4568,
    new_n4569, new_n4570, new_n4571, new_n4572, new_n4573, new_n4574,
    new_n4575, new_n4576, new_n4577, new_n4578, new_n4579, new_n4580,
    new_n4581, new_n4582, new_n4583, new_n4584, new_n4585, new_n4586,
    new_n4587, new_n4588, new_n4589, new_n4590, new_n4591, new_n4592,
    new_n4593, new_n4594, new_n4595, new_n4596, new_n4597, new_n4598,
    new_n4599, new_n4600, new_n4601, new_n4602, new_n4603, new_n4604,
    new_n4605, new_n4606, new_n4607, new_n4608, new_n4609, new_n4610,
    new_n4611, new_n4612, new_n4613, new_n4614, new_n4615, new_n4616,
    new_n4617, new_n4618, new_n4619, new_n4620, new_n4621, new_n4622,
    new_n4623, new_n4624, new_n4625, new_n4626, new_n4627, new_n4628,
    new_n4629, new_n4630, new_n4631, new_n4632, new_n4633, new_n4634,
    new_n4635, new_n4636, new_n4637, new_n4638, new_n4639, new_n4640,
    new_n4641, new_n4642, new_n4643, new_n4644, new_n4645, new_n4647,
    new_n4648, new_n4649, new_n4650, new_n4651, new_n4652, new_n4653,
    new_n4654, new_n4655, new_n4656, new_n4657, new_n4658, new_n4659,
    new_n4660, new_n4661, new_n4662, new_n4663, new_n4664, new_n4665,
    new_n4666, new_n4667, new_n4668, new_n4669, new_n4670, new_n4671,
    new_n4672, new_n4673, new_n4674, new_n4675, new_n4676, new_n4677,
    new_n4678, new_n4679, new_n4680, new_n4681, new_n4682, new_n4683,
    new_n4684, new_n4685, new_n4686, new_n4687, new_n4688, new_n4689,
    new_n4690, new_n4691, new_n4692, new_n4693, new_n4694, new_n4695,
    new_n4696, new_n4697, new_n4698, new_n4699, new_n4700, new_n4701,
    new_n4702, new_n4703, new_n4704, new_n4705, new_n4706, new_n4707,
    new_n4708, new_n4709, new_n4710, new_n4711, new_n4712, new_n4713,
    new_n4714, new_n4715, new_n4716, new_n4717, new_n4718, new_n4719,
    new_n4720, new_n4721, new_n4722, new_n4723, new_n4724, new_n4725,
    new_n4726, new_n4727, new_n4728, new_n4729, new_n4730, new_n4731,
    new_n4732, new_n4733, new_n4734, new_n4735, new_n4736, new_n4737,
    new_n4738, new_n4739, new_n4740, new_n4741, new_n4742, new_n4743,
    new_n4744, new_n4745, new_n4746, new_n4747, new_n4748, new_n4749,
    new_n4750, new_n4751, new_n4752, new_n4753, new_n4754, new_n4755,
    new_n4756, new_n4757, new_n4758, new_n4759, new_n4760, new_n4761,
    new_n4762, new_n4763, new_n4764, new_n4765, new_n4766, new_n4767,
    new_n4768, new_n4769, new_n4770, new_n4771, new_n4772, new_n4773,
    new_n4774, new_n4775, new_n4776, new_n4777, new_n4778, new_n4779,
    new_n4780, new_n4781, new_n4782, new_n4783, new_n4784, new_n4785,
    new_n4786, new_n4787, new_n4788, new_n4789, new_n4790, new_n4791,
    new_n4792, new_n4793, new_n4794, new_n4795, new_n4796, new_n4797,
    new_n4798, new_n4799, new_n4800, new_n4801, new_n4802, new_n4803,
    new_n4804, new_n4805, new_n4806, new_n4807, new_n4808, new_n4809,
    new_n4810, new_n4811, new_n4812, new_n4813, new_n4814, new_n4815,
    new_n4816, new_n4817, new_n4818, new_n4819, new_n4820, new_n4821,
    new_n4822, new_n4823, new_n4824, new_n4825, new_n4826, new_n4827,
    new_n4828, new_n4829, new_n4830, new_n4831, new_n4832, new_n4833,
    new_n4834, new_n4835, new_n4836, new_n4837, new_n4838, new_n4839,
    new_n4840, new_n4841, new_n4842, new_n4843, new_n4844, new_n4845,
    new_n4846, new_n4847, new_n4848, new_n4849, new_n4850, new_n4851,
    new_n4852, new_n4853, new_n4854, new_n4855, new_n4856, new_n4857,
    new_n4858, new_n4859, new_n4860, new_n4861, new_n4862, new_n4863,
    new_n4864, new_n4865, new_n4866, new_n4867, new_n4868, new_n4869,
    new_n4870, new_n4871, new_n4872, new_n4873, new_n4874, new_n4875,
    new_n4876, new_n4878, new_n4879, new_n4880, new_n4881, new_n4882,
    new_n4883, new_n4884, new_n4885, new_n4886, new_n4887, new_n4888,
    new_n4889, new_n4890, new_n4891, new_n4892, new_n4893, new_n4894,
    new_n4895, new_n4896, new_n4897, new_n4898, new_n4899, new_n4900,
    new_n4901, new_n4902, new_n4903, new_n4904, new_n4905, new_n4906,
    new_n4907, new_n4908, new_n4909, new_n4910, new_n4911, new_n4912,
    new_n4913, new_n4914, new_n4915, new_n4916, new_n4917, new_n4918,
    new_n4919, new_n4920, new_n4921, new_n4922, new_n4923, new_n4924,
    new_n4925, new_n4926, new_n4927, new_n4928, new_n4929, new_n4930,
    new_n4931, new_n4932, new_n4933, new_n4934, new_n4935, new_n4936,
    new_n4937, new_n4938, new_n4939, new_n4940, new_n4941, new_n4942,
    new_n4943, new_n4944, new_n4945, new_n4946, new_n4947, new_n4948,
    new_n4949, new_n4950, new_n4951, new_n4952, new_n4953, new_n4954,
    new_n4955, new_n4956, new_n4957, new_n4958, new_n4959, new_n4960,
    new_n4961, new_n4962, new_n4963, new_n4964, new_n4965, new_n4966,
    new_n4967, new_n4968, new_n4969, new_n4970, new_n4971, new_n4972,
    new_n4973, new_n4974, new_n4975, new_n4976, new_n4977, new_n4978,
    new_n4979, new_n4980, new_n4981, new_n4982, new_n4983, new_n4984,
    new_n4985, new_n4986, new_n4987, new_n4988, new_n4989, new_n4990,
    new_n4991, new_n4992, new_n4993, new_n4994, new_n4995, new_n4996,
    new_n4997, new_n4998, new_n4999, new_n5000, new_n5001, new_n5002,
    new_n5003, new_n5004, new_n5005, new_n5006, new_n5007, new_n5008,
    new_n5009, new_n5010, new_n5011, new_n5012, new_n5013, new_n5014,
    new_n5015, new_n5016, new_n5017, new_n5018, new_n5019, new_n5020,
    new_n5021, new_n5022, new_n5023, new_n5024, new_n5025, new_n5026,
    new_n5027, new_n5028, new_n5029, new_n5030, new_n5031, new_n5032,
    new_n5033, new_n5034, new_n5035, new_n5036, new_n5037, new_n5038,
    new_n5039, new_n5040, new_n5041, new_n5042, new_n5043, new_n5044,
    new_n5045, new_n5046, new_n5047, new_n5048, new_n5049, new_n5050,
    new_n5051, new_n5052, new_n5053, new_n5054, new_n5055, new_n5056,
    new_n5057, new_n5058, new_n5059, new_n5060, new_n5061, new_n5062,
    new_n5063, new_n5064, new_n5065, new_n5066, new_n5067, new_n5068,
    new_n5069, new_n5070, new_n5071, new_n5072, new_n5073, new_n5074,
    new_n5075, new_n5076, new_n5077, new_n5078, new_n5079, new_n5080,
    new_n5081, new_n5082, new_n5083, new_n5084, new_n5085, new_n5086,
    new_n5087, new_n5088, new_n5089, new_n5090, new_n5091, new_n5092,
    new_n5093, new_n5094, new_n5095, new_n5096, new_n5097, new_n5098,
    new_n5099, new_n5100, new_n5101, new_n5102, new_n5103, new_n5104,
    new_n5105, new_n5106, new_n5107, new_n5108, new_n5109, new_n5110,
    new_n5111, new_n5112, new_n5113, new_n5114, new_n5115, new_n5116,
    new_n5117, new_n5118, new_n5119, new_n5121, new_n5122, new_n5123,
    new_n5124, new_n5125, new_n5126, new_n5127, new_n5128, new_n5129,
    new_n5130, new_n5131, new_n5132, new_n5133, new_n5134, new_n5135,
    new_n5136, new_n5137, new_n5138, new_n5139, new_n5140, new_n5141,
    new_n5142, new_n5143, new_n5144, new_n5145, new_n5146, new_n5147,
    new_n5148, new_n5149, new_n5150, new_n5151, new_n5152, new_n5153,
    new_n5154, new_n5155, new_n5156, new_n5157, new_n5158, new_n5159,
    new_n5160, new_n5161, new_n5162, new_n5163, new_n5164, new_n5165,
    new_n5166, new_n5167, new_n5168, new_n5169, new_n5170, new_n5171,
    new_n5172, new_n5173, new_n5174, new_n5175, new_n5176, new_n5177,
    new_n5178, new_n5179, new_n5180, new_n5181, new_n5182, new_n5183,
    new_n5184, new_n5185, new_n5186, new_n5187, new_n5188, new_n5189,
    new_n5190, new_n5191, new_n5192, new_n5193, new_n5194, new_n5195,
    new_n5196, new_n5197, new_n5198, new_n5199, new_n5200, new_n5201,
    new_n5202, new_n5203, new_n5204, new_n5205, new_n5206, new_n5207,
    new_n5208, new_n5209, new_n5210, new_n5211, new_n5212, new_n5213,
    new_n5214, new_n5215, new_n5216, new_n5217, new_n5218, new_n5219,
    new_n5220, new_n5221, new_n5222, new_n5223, new_n5224, new_n5225,
    new_n5226, new_n5227, new_n5228, new_n5229, new_n5230, new_n5231,
    new_n5232, new_n5233, new_n5234, new_n5235, new_n5236, new_n5237,
    new_n5238, new_n5239, new_n5240, new_n5241, new_n5242, new_n5243,
    new_n5244, new_n5245, new_n5246, new_n5247, new_n5248, new_n5249,
    new_n5250, new_n5251, new_n5252, new_n5253, new_n5254, new_n5255,
    new_n5256, new_n5257, new_n5258, new_n5259, new_n5260, new_n5261,
    new_n5262, new_n5263, new_n5264, new_n5265, new_n5266, new_n5267,
    new_n5268, new_n5269, new_n5270, new_n5271, new_n5272, new_n5273,
    new_n5274, new_n5275, new_n5276, new_n5277, new_n5278, new_n5279,
    new_n5280, new_n5281, new_n5282, new_n5283, new_n5284, new_n5285,
    new_n5286, new_n5287, new_n5288, new_n5289, new_n5290, new_n5291,
    new_n5292, new_n5293, new_n5294, new_n5295, new_n5296, new_n5297,
    new_n5298, new_n5299, new_n5300, new_n5301, new_n5302, new_n5303,
    new_n5304, new_n5305, new_n5306, new_n5307, new_n5308, new_n5309,
    new_n5310, new_n5311, new_n5312, new_n5313, new_n5314, new_n5315,
    new_n5316, new_n5317, new_n5318, new_n5319, new_n5320, new_n5321,
    new_n5322, new_n5323, new_n5324, new_n5325, new_n5326, new_n5327,
    new_n5328, new_n5329, new_n5330, new_n5331, new_n5332, new_n5333,
    new_n5334, new_n5335, new_n5336, new_n5337, new_n5338, new_n5339,
    new_n5340, new_n5341, new_n5342, new_n5343, new_n5344, new_n5345,
    new_n5346, new_n5347, new_n5348, new_n5349, new_n5350, new_n5351,
    new_n5352, new_n5353, new_n5354, new_n5355, new_n5356, new_n5357,
    new_n5358, new_n5359, new_n5360, new_n5361, new_n5363, new_n5364,
    new_n5365, new_n5366, new_n5367, new_n5368, new_n5369, new_n5370,
    new_n5371, new_n5372, new_n5373, new_n5374, new_n5375, new_n5376,
    new_n5377, new_n5378, new_n5379, new_n5380, new_n5381, new_n5382,
    new_n5383, new_n5384, new_n5385, new_n5386, new_n5387, new_n5388,
    new_n5389, new_n5390, new_n5391, new_n5392, new_n5393, new_n5394,
    new_n5395, new_n5396, new_n5397, new_n5398, new_n5399, new_n5400,
    new_n5401, new_n5402, new_n5403, new_n5404, new_n5405, new_n5406,
    new_n5407, new_n5408, new_n5409, new_n5410, new_n5411, new_n5412,
    new_n5413, new_n5414, new_n5415, new_n5416, new_n5417, new_n5418,
    new_n5419, new_n5420, new_n5421, new_n5422, new_n5423, new_n5424,
    new_n5425, new_n5426, new_n5427, new_n5428, new_n5429, new_n5430,
    new_n5431, new_n5432, new_n5433, new_n5434, new_n5435, new_n5436,
    new_n5437, new_n5438, new_n5439, new_n5440, new_n5441, new_n5442,
    new_n5443, new_n5444, new_n5445, new_n5446, new_n5447, new_n5448,
    new_n5449, new_n5450, new_n5451, new_n5452, new_n5453, new_n5454,
    new_n5455, new_n5456, new_n5457, new_n5458, new_n5459, new_n5460,
    new_n5461, new_n5462, new_n5463, new_n5464, new_n5465, new_n5466,
    new_n5467, new_n5468, new_n5469, new_n5470, new_n5471, new_n5472,
    new_n5473, new_n5474, new_n5475, new_n5476, new_n5477, new_n5478,
    new_n5479, new_n5480, new_n5481, new_n5482, new_n5483, new_n5484,
    new_n5485, new_n5486, new_n5487, new_n5488, new_n5489, new_n5490,
    new_n5491, new_n5492, new_n5493, new_n5494, new_n5495, new_n5496,
    new_n5497, new_n5498, new_n5499, new_n5500, new_n5501, new_n5502,
    new_n5503, new_n5504, new_n5505, new_n5506, new_n5507, new_n5508,
    new_n5509, new_n5510, new_n5511, new_n5512, new_n5513, new_n5514,
    new_n5515, new_n5516, new_n5517, new_n5518, new_n5519, new_n5520,
    new_n5521, new_n5522, new_n5523, new_n5524, new_n5525, new_n5526,
    new_n5527, new_n5528, new_n5529, new_n5530, new_n5531, new_n5532,
    new_n5533, new_n5534, new_n5535, new_n5536, new_n5537, new_n5538,
    new_n5539, new_n5540, new_n5541, new_n5542, new_n5543, new_n5544,
    new_n5545, new_n5546, new_n5547, new_n5548, new_n5549, new_n5550,
    new_n5551, new_n5552, new_n5553, new_n5554, new_n5555, new_n5556,
    new_n5557, new_n5558, new_n5559, new_n5560, new_n5561, new_n5562,
    new_n5563, new_n5564, new_n5565, new_n5566, new_n5567, new_n5568,
    new_n5569, new_n5570, new_n5571, new_n5572, new_n5573, new_n5574,
    new_n5575, new_n5576, new_n5577, new_n5578, new_n5579, new_n5580,
    new_n5581, new_n5582, new_n5583, new_n5584, new_n5585, new_n5586,
    new_n5587, new_n5588, new_n5589, new_n5590, new_n5591, new_n5592,
    new_n5593, new_n5594, new_n5595, new_n5596, new_n5597, new_n5598,
    new_n5599, new_n5600, new_n5601, new_n5602, new_n5603, new_n5604,
    new_n5605, new_n5606, new_n5607, new_n5608, new_n5609, new_n5610,
    new_n5611, new_n5613, new_n5614, new_n5615, new_n5616, new_n5617,
    new_n5618, new_n5619, new_n5620, new_n5621, new_n5622, new_n5623,
    new_n5624, new_n5625, new_n5626, new_n5627, new_n5628, new_n5629,
    new_n5630, new_n5631, new_n5632, new_n5633, new_n5634, new_n5635,
    new_n5636, new_n5637, new_n5638, new_n5639, new_n5640, new_n5641,
    new_n5642, new_n5643, new_n5644, new_n5645, new_n5646, new_n5647,
    new_n5648, new_n5649, new_n5650, new_n5651, new_n5652, new_n5653,
    new_n5654, new_n5655, new_n5656, new_n5657, new_n5658, new_n5659,
    new_n5660, new_n5661, new_n5662, new_n5663, new_n5664, new_n5665,
    new_n5666, new_n5667, new_n5668, new_n5669, new_n5670, new_n5671,
    new_n5672, new_n5673, new_n5674, new_n5675, new_n5676, new_n5677,
    new_n5678, new_n5679, new_n5680, new_n5681, new_n5682, new_n5683,
    new_n5684, new_n5685, new_n5686, new_n5687, new_n5688, new_n5689,
    new_n5690, new_n5691, new_n5692, new_n5693, new_n5694, new_n5695,
    new_n5696, new_n5697, new_n5698, new_n5699, new_n5700, new_n5701,
    new_n5702, new_n5703, new_n5704, new_n5705, new_n5706, new_n5707,
    new_n5708, new_n5709, new_n5710, new_n5711, new_n5712, new_n5713,
    new_n5714, new_n5715, new_n5716, new_n5717, new_n5718, new_n5719,
    new_n5720, new_n5721, new_n5722, new_n5723, new_n5724, new_n5725,
    new_n5726, new_n5727, new_n5728, new_n5729, new_n5730, new_n5731,
    new_n5732, new_n5733, new_n5734, new_n5735, new_n5736, new_n5737,
    new_n5738, new_n5739, new_n5740, new_n5741, new_n5742, new_n5743,
    new_n5744, new_n5745, new_n5746, new_n5747, new_n5748, new_n5749,
    new_n5750, new_n5751, new_n5752, new_n5753, new_n5754, new_n5755,
    new_n5756, new_n5757, new_n5758, new_n5759, new_n5760, new_n5761,
    new_n5762, new_n5763, new_n5764, new_n5765, new_n5766, new_n5767,
    new_n5768, new_n5769, new_n5770, new_n5771, new_n5772, new_n5773,
    new_n5774, new_n5775, new_n5776, new_n5777, new_n5778, new_n5779,
    new_n5780, new_n5781, new_n5782, new_n5783, new_n5784, new_n5785,
    new_n5786, new_n5787, new_n5788, new_n5789, new_n5790, new_n5791,
    new_n5792, new_n5793, new_n5794, new_n5795, new_n5796, new_n5797,
    new_n5798, new_n5799, new_n5800, new_n5801, new_n5802, new_n5803,
    new_n5804, new_n5805, new_n5806, new_n5807, new_n5808, new_n5809,
    new_n5810, new_n5811, new_n5812, new_n5813, new_n5814, new_n5815,
    new_n5816, new_n5817, new_n5818, new_n5819, new_n5820, new_n5821,
    new_n5822, new_n5823, new_n5824, new_n5825, new_n5826, new_n5827,
    new_n5828, new_n5829, new_n5830, new_n5831, new_n5832, new_n5833,
    new_n5834, new_n5835, new_n5836, new_n5837, new_n5838, new_n5839,
    new_n5840, new_n5841, new_n5842, new_n5843, new_n5844, new_n5845,
    new_n5846, new_n5847, new_n5848, new_n5849, new_n5850, new_n5851,
    new_n5852, new_n5853, new_n5854, new_n5855, new_n5856, new_n5857,
    new_n5858, new_n5859, new_n5860, new_n5861, new_n5862, new_n5864,
    new_n5865, new_n5866, new_n5867, new_n5868, new_n5869, new_n5870,
    new_n5871, new_n5872, new_n5873, new_n5874, new_n5875, new_n5876,
    new_n5877, new_n5878, new_n5879, new_n5880, new_n5881, new_n5882,
    new_n5883, new_n5884, new_n5885, new_n5886, new_n5887, new_n5888,
    new_n5889, new_n5890, new_n5891, new_n5892, new_n5893, new_n5894,
    new_n5895, new_n5896, new_n5897, new_n5898, new_n5899, new_n5900,
    new_n5901, new_n5902, new_n5903, new_n5904, new_n5905, new_n5906,
    new_n5907, new_n5908, new_n5909, new_n5910, new_n5911, new_n5912,
    new_n5913, new_n5914, new_n5915, new_n5916, new_n5917, new_n5918,
    new_n5919, new_n5920, new_n5921, new_n5922, new_n5923, new_n5924,
    new_n5925, new_n5926, new_n5927, new_n5928, new_n5929, new_n5930,
    new_n5931, new_n5932, new_n5933, new_n5934, new_n5935, new_n5936,
    new_n5937, new_n5938, new_n5939, new_n5940, new_n5941, new_n5942,
    new_n5943, new_n5944, new_n5945, new_n5946, new_n5947, new_n5948,
    new_n5949, new_n5950, new_n5951, new_n5952, new_n5953, new_n5954,
    new_n5955, new_n5956, new_n5957, new_n5958, new_n5959, new_n5960,
    new_n5961, new_n5962, new_n5963, new_n5964, new_n5965, new_n5966,
    new_n5967, new_n5968, new_n5969, new_n5970, new_n5971, new_n5972,
    new_n5973, new_n5974, new_n5975, new_n5976, new_n5977, new_n5978,
    new_n5979, new_n5980, new_n5981, new_n5982, new_n5983, new_n5984,
    new_n5985, new_n5986, new_n5987, new_n5988, new_n5989, new_n5990,
    new_n5991, new_n5992, new_n5993, new_n5994, new_n5995, new_n5996,
    new_n5997, new_n5998, new_n5999, new_n6000, new_n6001, new_n6002,
    new_n6003, new_n6004, new_n6005, new_n6006, new_n6007, new_n6008,
    new_n6009, new_n6010, new_n6011, new_n6012, new_n6013, new_n6014,
    new_n6015, new_n6016, new_n6017, new_n6018, new_n6019, new_n6020,
    new_n6021, new_n6022, new_n6023, new_n6024, new_n6025, new_n6026,
    new_n6027, new_n6028, new_n6029, new_n6030, new_n6031, new_n6032,
    new_n6033, new_n6034, new_n6035, new_n6036, new_n6037, new_n6038,
    new_n6039, new_n6040, new_n6041, new_n6042, new_n6043, new_n6044,
    new_n6045, new_n6046, new_n6047, new_n6048, new_n6049, new_n6050,
    new_n6051, new_n6052, new_n6053, new_n6054, new_n6055, new_n6056,
    new_n6057, new_n6058, new_n6059, new_n6060, new_n6061, new_n6062,
    new_n6063, new_n6064, new_n6065, new_n6066, new_n6067, new_n6068,
    new_n6069, new_n6070, new_n6071, new_n6072, new_n6073, new_n6074,
    new_n6075, new_n6076, new_n6077, new_n6078, new_n6079, new_n6080,
    new_n6081, new_n6082, new_n6083, new_n6084, new_n6085, new_n6086,
    new_n6087, new_n6088, new_n6089, new_n6090, new_n6091, new_n6092,
    new_n6093, new_n6094, new_n6095, new_n6096, new_n6097, new_n6098,
    new_n6099, new_n6100, new_n6101, new_n6102, new_n6103, new_n6104,
    new_n6105, new_n6106, new_n6107, new_n6108, new_n6109, new_n6110,
    new_n6111, new_n6112, new_n6113, new_n6114, new_n6115, new_n6116,
    new_n6117, new_n6118, new_n6119, new_n6120, new_n6121, new_n6122,
    new_n6123, new_n6125, new_n6126, new_n6127, new_n6128, new_n6129,
    new_n6130, new_n6131, new_n6132, new_n6133, new_n6134, new_n6135,
    new_n6136, new_n6137, new_n6138, new_n6139, new_n6140, new_n6141,
    new_n6142, new_n6143, new_n6144, new_n6145, new_n6146, new_n6147,
    new_n6148, new_n6149, new_n6150, new_n6151, new_n6152, new_n6153,
    new_n6154, new_n6155, new_n6156, new_n6157, new_n6158, new_n6159,
    new_n6160, new_n6161, new_n6162, new_n6163, new_n6164, new_n6165,
    new_n6166, new_n6167, new_n6168, new_n6169, new_n6170, new_n6171,
    new_n6172, new_n6173, new_n6174, new_n6175, new_n6176, new_n6177,
    new_n6178, new_n6179, new_n6180, new_n6181, new_n6182, new_n6183,
    new_n6184, new_n6185, new_n6186, new_n6187, new_n6188, new_n6189,
    new_n6190, new_n6191, new_n6192, new_n6193, new_n6194, new_n6195,
    new_n6196, new_n6197, new_n6198, new_n6199, new_n6200, new_n6201,
    new_n6202, new_n6203, new_n6204, new_n6205, new_n6206, new_n6207,
    new_n6208, new_n6209, new_n6210, new_n6211, new_n6212, new_n6213,
    new_n6214, new_n6215, new_n6216, new_n6217, new_n6218, new_n6219,
    new_n6220, new_n6221, new_n6222, new_n6223, new_n6224, new_n6225,
    new_n6226, new_n6227, new_n6228, new_n6229, new_n6230, new_n6231,
    new_n6232, new_n6233, new_n6234, new_n6235, new_n6236, new_n6237,
    new_n6238, new_n6239, new_n6240, new_n6241, new_n6242, new_n6243,
    new_n6244, new_n6245, new_n6246, new_n6247, new_n6248, new_n6249,
    new_n6250, new_n6251, new_n6252, new_n6253, new_n6254, new_n6255,
    new_n6256, new_n6257, new_n6258, new_n6259, new_n6260, new_n6261,
    new_n6262, new_n6263, new_n6264, new_n6265, new_n6266, new_n6267,
    new_n6268, new_n6269, new_n6270, new_n6271, new_n6272, new_n6273,
    new_n6274, new_n6275, new_n6276, new_n6277, new_n6278, new_n6279,
    new_n6280, new_n6281, new_n6282, new_n6283, new_n6284, new_n6285,
    new_n6286, new_n6287, new_n6288, new_n6289, new_n6290, new_n6291,
    new_n6292, new_n6293, new_n6294, new_n6295, new_n6296, new_n6297,
    new_n6298, new_n6299, new_n6300, new_n6301, new_n6302, new_n6303,
    new_n6304, new_n6305, new_n6306, new_n6307, new_n6308, new_n6309,
    new_n6310, new_n6311, new_n6312, new_n6313, new_n6314, new_n6315,
    new_n6316, new_n6317, new_n6318, new_n6319, new_n6320, new_n6321,
    new_n6322, new_n6323, new_n6324, new_n6325, new_n6326, new_n6327,
    new_n6328, new_n6329, new_n6330, new_n6331, new_n6332, new_n6333,
    new_n6334, new_n6335, new_n6336, new_n6337, new_n6338, new_n6339,
    new_n6340, new_n6341, new_n6342, new_n6343, new_n6344, new_n6345,
    new_n6346, new_n6347, new_n6348, new_n6349, new_n6350, new_n6351,
    new_n6352, new_n6353, new_n6354, new_n6355, new_n6356, new_n6357,
    new_n6358, new_n6359, new_n6360, new_n6361, new_n6362, new_n6363,
    new_n6364, new_n6365, new_n6366, new_n6367, new_n6368, new_n6369,
    new_n6370, new_n6371, new_n6372, new_n6373, new_n6374, new_n6375,
    new_n6376, new_n6377, new_n6378, new_n6379, new_n6380, new_n6381,
    new_n6382, new_n6383, new_n6384, new_n6385, new_n6386, new_n6387,
    new_n6388, new_n6390, new_n6391, new_n6392, new_n6393, new_n6394,
    new_n6395, new_n6396, new_n6397, new_n6398, new_n6399, new_n6400,
    new_n6401, new_n6402, new_n6403, new_n6404, new_n6405, new_n6406,
    new_n6407, new_n6408, new_n6409, new_n6410, new_n6411, new_n6412,
    new_n6413, new_n6414, new_n6415, new_n6416, new_n6417, new_n6418,
    new_n6419, new_n6420, new_n6421, new_n6422, new_n6423, new_n6424,
    new_n6425, new_n6426, new_n6427, new_n6428, new_n6429, new_n6430,
    new_n6431, new_n6432, new_n6433, new_n6434, new_n6435, new_n6436,
    new_n6437, new_n6438, new_n6439, new_n6440, new_n6441, new_n6442,
    new_n6443, new_n6444, new_n6445, new_n6446, new_n6447, new_n6448,
    new_n6449, new_n6450, new_n6451, new_n6452, new_n6453, new_n6454,
    new_n6455, new_n6456, new_n6457, new_n6458, new_n6459, new_n6460,
    new_n6461, new_n6462, new_n6463, new_n6464, new_n6465, new_n6466,
    new_n6467, new_n6468, new_n6469, new_n6470, new_n6471, new_n6472,
    new_n6473, new_n6474, new_n6475, new_n6476, new_n6477, new_n6478,
    new_n6479, new_n6480, new_n6481, new_n6482, new_n6483, new_n6484,
    new_n6485, new_n6486, new_n6487, new_n6488, new_n6489, new_n6490,
    new_n6491, new_n6492, new_n6493, new_n6494, new_n6495, new_n6496,
    new_n6497, new_n6498, new_n6499, new_n6500, new_n6501, new_n6502,
    new_n6503, new_n6504, new_n6505, new_n6506, new_n6507, new_n6508,
    new_n6509, new_n6510, new_n6511, new_n6512, new_n6513, new_n6514,
    new_n6515, new_n6516, new_n6517, new_n6518, new_n6519, new_n6520,
    new_n6521, new_n6522, new_n6523, new_n6524, new_n6525, new_n6526,
    new_n6527, new_n6528, new_n6529, new_n6530, new_n6531, new_n6532,
    new_n6533, new_n6534, new_n6535, new_n6536, new_n6537, new_n6538,
    new_n6539, new_n6540, new_n6541, new_n6542, new_n6543, new_n6544,
    new_n6545, new_n6546, new_n6547, new_n6548, new_n6549, new_n6550,
    new_n6551, new_n6552, new_n6553, new_n6554, new_n6555, new_n6556,
    new_n6557, new_n6558, new_n6559, new_n6560, new_n6561, new_n6562,
    new_n6563, new_n6564, new_n6565, new_n6566, new_n6567, new_n6568,
    new_n6569, new_n6570, new_n6571, new_n6572, new_n6573, new_n6574,
    new_n6575, new_n6576, new_n6577, new_n6578, new_n6579, new_n6580,
    new_n6581, new_n6582, new_n6583, new_n6584, new_n6585, new_n6586,
    new_n6587, new_n6588, new_n6589, new_n6590, new_n6591, new_n6592,
    new_n6593, new_n6594, new_n6595, new_n6596, new_n6597, new_n6598,
    new_n6599, new_n6600, new_n6601, new_n6602, new_n6603, new_n6604,
    new_n6605, new_n6606, new_n6607, new_n6608, new_n6609, new_n6610,
    new_n6611, new_n6612, new_n6613, new_n6614, new_n6615, new_n6616,
    new_n6617, new_n6618, new_n6619, new_n6620, new_n6621, new_n6622,
    new_n6623, new_n6624, new_n6625, new_n6626, new_n6627, new_n6628,
    new_n6629, new_n6630, new_n6631, new_n6632, new_n6633, new_n6634,
    new_n6635, new_n6636, new_n6637, new_n6638, new_n6639, new_n6640,
    new_n6641, new_n6642, new_n6643, new_n6644, new_n6645, new_n6646,
    new_n6647, new_n6648, new_n6649, new_n6650, new_n6651, new_n6652,
    new_n6653, new_n6654, new_n6655, new_n6656, new_n6657, new_n6658,
    new_n6659, new_n6660, new_n6661, new_n6662, new_n6663, new_n6664,
    new_n6665, new_n6666, new_n6668, new_n6669, new_n6670, new_n6671,
    new_n6672, new_n6673, new_n6674, new_n6675, new_n6676, new_n6677,
    new_n6678, new_n6679, new_n6680, new_n6681, new_n6682, new_n6683,
    new_n6684, new_n6685, new_n6686, new_n6687, new_n6688, new_n6689,
    new_n6690, new_n6691, new_n6692, new_n6693, new_n6694, new_n6695,
    new_n6696, new_n6697, new_n6698, new_n6699, new_n6700, new_n6701,
    new_n6702, new_n6703, new_n6704, new_n6705, new_n6706, new_n6707,
    new_n6708, new_n6709, new_n6710, new_n6711, new_n6712, new_n6713,
    new_n6714, new_n6715, new_n6716, new_n6717, new_n6718, new_n6719,
    new_n6720, new_n6721, new_n6722, new_n6723, new_n6724, new_n6725,
    new_n6726, new_n6727, new_n6728, new_n6729, new_n6730, new_n6731,
    new_n6732, new_n6733, new_n6734, new_n6735, new_n6736, new_n6737,
    new_n6738, new_n6739, new_n6740, new_n6741, new_n6742, new_n6743,
    new_n6744, new_n6745, new_n6746, new_n6747, new_n6748, new_n6749,
    new_n6750, new_n6751, new_n6752, new_n6753, new_n6754, new_n6755,
    new_n6756, new_n6757, new_n6758, new_n6759, new_n6760, new_n6761,
    new_n6762, new_n6763, new_n6764, new_n6765, new_n6766, new_n6767,
    new_n6768, new_n6769, new_n6770, new_n6771, new_n6772, new_n6773,
    new_n6774, new_n6775, new_n6776, new_n6777, new_n6778, new_n6779,
    new_n6780, new_n6781, new_n6782, new_n6783, new_n6784, new_n6785,
    new_n6786, new_n6787, new_n6788, new_n6789, new_n6790, new_n6791,
    new_n6792, new_n6793, new_n6794, new_n6795, new_n6796, new_n6797,
    new_n6798, new_n6799, new_n6800, new_n6801, new_n6802, new_n6803,
    new_n6804, new_n6805, new_n6806, new_n6807, new_n6808, new_n6809,
    new_n6810, new_n6811, new_n6812, new_n6813, new_n6814, new_n6815,
    new_n6816, new_n6817, new_n6818, new_n6819, new_n6820, new_n6821,
    new_n6822, new_n6823, new_n6824, new_n6825, new_n6826, new_n6827,
    new_n6828, new_n6829, new_n6830, new_n6831, new_n6832, new_n6833,
    new_n6834, new_n6835, new_n6836, new_n6837, new_n6838, new_n6839,
    new_n6840, new_n6841, new_n6842, new_n6843, new_n6844, new_n6845,
    new_n6846, new_n6847, new_n6848, new_n6849, new_n6850, new_n6851,
    new_n6852, new_n6853, new_n6854, new_n6855, new_n6856, new_n6857,
    new_n6858, new_n6859, new_n6860, new_n6861, new_n6862, new_n6863,
    new_n6864, new_n6865, new_n6866, new_n6867, new_n6868, new_n6869,
    new_n6870, new_n6871, new_n6872, new_n6873, new_n6874, new_n6875,
    new_n6876, new_n6877, new_n6878, new_n6879, new_n6880, new_n6881,
    new_n6882, new_n6883, new_n6884, new_n6885, new_n6886, new_n6887,
    new_n6888, new_n6889, new_n6890, new_n6891, new_n6892, new_n6893,
    new_n6894, new_n6895, new_n6896, new_n6897, new_n6898, new_n6899,
    new_n6900, new_n6901, new_n6902, new_n6903, new_n6904, new_n6905,
    new_n6906, new_n6907, new_n6908, new_n6909, new_n6910, new_n6911,
    new_n6912, new_n6913, new_n6914, new_n6915, new_n6916, new_n6917,
    new_n6918, new_n6919, new_n6920, new_n6921, new_n6922, new_n6923,
    new_n6924, new_n6925, new_n6926, new_n6927, new_n6928, new_n6929,
    new_n6930, new_n6931, new_n6932, new_n6933, new_n6934, new_n6935,
    new_n6936, new_n6937, new_n6938, new_n6939, new_n6941, new_n6942,
    new_n6943, new_n6944, new_n6945, new_n6946, new_n6947, new_n6948,
    new_n6949, new_n6950, new_n6951, new_n6952, new_n6953, new_n6954,
    new_n6955, new_n6956, new_n6957, new_n6958, new_n6959, new_n6960,
    new_n6961, new_n6962, new_n6963, new_n6964, new_n6965, new_n6966,
    new_n6967, new_n6968, new_n6969, new_n6970, new_n6971, new_n6972,
    new_n6973, new_n6974, new_n6975, new_n6976, new_n6977, new_n6978,
    new_n6979, new_n6980, new_n6981, new_n6982, new_n6983, new_n6984,
    new_n6985, new_n6986, new_n6987, new_n6988, new_n6989, new_n6990,
    new_n6991, new_n6992, new_n6993, new_n6994, new_n6995, new_n6996,
    new_n6997, new_n6998, new_n6999, new_n7000, new_n7001, new_n7002,
    new_n7003, new_n7004, new_n7005, new_n7006, new_n7007, new_n7008,
    new_n7009, new_n7010, new_n7011, new_n7012, new_n7013, new_n7014,
    new_n7015, new_n7016, new_n7017, new_n7018, new_n7019, new_n7020,
    new_n7021, new_n7022, new_n7023, new_n7024, new_n7025, new_n7026,
    new_n7027, new_n7028, new_n7029, new_n7030, new_n7031, new_n7032,
    new_n7033, new_n7034, new_n7035, new_n7036, new_n7037, new_n7038,
    new_n7039, new_n7040, new_n7041, new_n7042, new_n7043, new_n7044,
    new_n7045, new_n7046, new_n7047, new_n7048, new_n7049, new_n7050,
    new_n7051, new_n7052, new_n7053, new_n7054, new_n7055, new_n7056,
    new_n7057, new_n7058, new_n7059, new_n7060, new_n7061, new_n7062,
    new_n7063, new_n7064, new_n7065, new_n7066, new_n7067, new_n7068,
    new_n7069, new_n7070, new_n7071, new_n7072, new_n7073, new_n7074,
    new_n7075, new_n7076, new_n7077, new_n7078, new_n7079, new_n7080,
    new_n7081, new_n7082, new_n7083, new_n7084, new_n7085, new_n7086,
    new_n7087, new_n7088, new_n7089, new_n7090, new_n7091, new_n7092,
    new_n7093, new_n7094, new_n7095, new_n7096, new_n7097, new_n7098,
    new_n7099, new_n7100, new_n7101, new_n7102, new_n7103, new_n7104,
    new_n7105, new_n7106, new_n7107, new_n7108, new_n7109, new_n7110,
    new_n7111, new_n7112, new_n7113, new_n7114, new_n7115, new_n7116,
    new_n7117, new_n7118, new_n7119, new_n7120, new_n7121, new_n7122,
    new_n7123, new_n7124, new_n7125, new_n7126, new_n7127, new_n7128,
    new_n7129, new_n7130, new_n7131, new_n7132, new_n7133, new_n7134,
    new_n7135, new_n7136, new_n7137, new_n7138, new_n7139, new_n7140,
    new_n7141, new_n7142, new_n7143, new_n7144, new_n7145, new_n7146,
    new_n7147, new_n7148, new_n7149, new_n7150, new_n7151, new_n7152,
    new_n7153, new_n7154, new_n7155, new_n7156, new_n7157, new_n7158,
    new_n7159, new_n7160, new_n7161, new_n7162, new_n7163, new_n7164,
    new_n7165, new_n7166, new_n7167, new_n7168, new_n7169, new_n7170,
    new_n7171, new_n7172, new_n7173, new_n7174, new_n7175, new_n7176,
    new_n7177, new_n7178, new_n7179, new_n7180, new_n7181, new_n7182,
    new_n7183, new_n7184, new_n7185, new_n7186, new_n7187, new_n7188,
    new_n7189, new_n7190, new_n7191, new_n7192, new_n7193, new_n7194,
    new_n7195, new_n7196, new_n7197, new_n7198, new_n7199, new_n7200,
    new_n7201, new_n7202, new_n7203, new_n7204, new_n7205, new_n7206,
    new_n7207, new_n7208, new_n7209, new_n7210, new_n7211, new_n7212,
    new_n7213, new_n7214, new_n7215, new_n7216, new_n7217, new_n7218,
    new_n7219, new_n7220, new_n7221, new_n7222, new_n7223, new_n7224,
    new_n7225, new_n7227, new_n7228, new_n7229, new_n7230, new_n7231,
    new_n7232, new_n7233, new_n7234, new_n7235, new_n7236, new_n7237,
    new_n7238, new_n7239, new_n7240, new_n7241, new_n7242, new_n7243,
    new_n7244, new_n7245, new_n7246, new_n7247, new_n7248, new_n7249,
    new_n7250, new_n7251, new_n7252, new_n7253, new_n7254, new_n7255,
    new_n7256, new_n7257, new_n7258, new_n7259, new_n7260, new_n7261,
    new_n7262, new_n7263, new_n7264, new_n7265, new_n7266, new_n7267,
    new_n7268, new_n7269, new_n7270, new_n7271, new_n7272, new_n7273,
    new_n7274, new_n7275, new_n7276, new_n7277, new_n7278, new_n7279,
    new_n7280, new_n7281, new_n7282, new_n7283, new_n7284, new_n7285,
    new_n7286, new_n7287, new_n7288, new_n7289, new_n7290, new_n7291,
    new_n7292, new_n7293, new_n7294, new_n7295, new_n7296, new_n7297,
    new_n7298, new_n7299, new_n7300, new_n7301, new_n7302, new_n7303,
    new_n7304, new_n7305, new_n7306, new_n7307, new_n7308, new_n7309,
    new_n7310, new_n7311, new_n7312, new_n7313, new_n7314, new_n7315,
    new_n7316, new_n7317, new_n7318, new_n7319, new_n7320, new_n7321,
    new_n7322, new_n7323, new_n7324, new_n7325, new_n7326, new_n7327,
    new_n7328, new_n7329, new_n7330, new_n7331, new_n7332, new_n7333,
    new_n7334, new_n7335, new_n7336, new_n7337, new_n7338, new_n7339,
    new_n7340, new_n7341, new_n7342, new_n7343, new_n7344, new_n7345,
    new_n7346, new_n7347, new_n7348, new_n7349, new_n7350, new_n7351,
    new_n7352, new_n7353, new_n7354, new_n7355, new_n7356, new_n7357,
    new_n7358, new_n7359, new_n7360, new_n7361, new_n7362, new_n7363,
    new_n7364, new_n7365, new_n7366, new_n7367, new_n7368, new_n7369,
    new_n7370, new_n7371, new_n7372, new_n7373, new_n7374, new_n7375,
    new_n7376, new_n7377, new_n7378, new_n7379, new_n7380, new_n7381,
    new_n7382, new_n7383, new_n7384, new_n7385, new_n7386, new_n7387,
    new_n7388, new_n7389, new_n7390, new_n7391, new_n7392, new_n7393,
    new_n7394, new_n7395, new_n7396, new_n7397, new_n7398, new_n7399,
    new_n7400, new_n7401, new_n7402, new_n7403, new_n7404, new_n7405,
    new_n7406, new_n7407, new_n7408, new_n7409, new_n7410, new_n7411,
    new_n7412, new_n7413, new_n7414, new_n7415, new_n7416, new_n7417,
    new_n7418, new_n7419, new_n7420, new_n7421, new_n7422, new_n7423,
    new_n7424, new_n7425, new_n7426, new_n7427, new_n7428, new_n7429,
    new_n7430, new_n7431, new_n7432, new_n7433, new_n7434, new_n7435,
    new_n7436, new_n7437, new_n7438, new_n7439, new_n7440, new_n7441,
    new_n7442, new_n7443, new_n7444, new_n7445, new_n7446, new_n7447,
    new_n7448, new_n7449, new_n7450, new_n7451, new_n7452, new_n7453,
    new_n7454, new_n7455, new_n7456, new_n7457, new_n7458, new_n7459,
    new_n7460, new_n7461, new_n7462, new_n7463, new_n7464, new_n7465,
    new_n7466, new_n7467, new_n7468, new_n7469, new_n7470, new_n7471,
    new_n7472, new_n7473, new_n7474, new_n7475, new_n7476, new_n7477,
    new_n7478, new_n7479, new_n7480, new_n7481, new_n7482, new_n7483,
    new_n7484, new_n7485, new_n7486, new_n7487, new_n7488, new_n7489,
    new_n7490, new_n7491, new_n7492, new_n7493, new_n7494, new_n7495,
    new_n7496, new_n7497, new_n7498, new_n7499, new_n7500, new_n7501,
    new_n7502, new_n7503, new_n7504, new_n7505, new_n7506, new_n7507,
    new_n7508, new_n7509, new_n7510, new_n7511, new_n7512, new_n7513,
    new_n7514, new_n7515, new_n7517, new_n7518, new_n7519, new_n7520,
    new_n7521, new_n7522, new_n7523, new_n7524, new_n7525, new_n7526,
    new_n7527, new_n7528, new_n7529, new_n7530, new_n7531, new_n7532,
    new_n7533, new_n7534, new_n7535, new_n7536, new_n7537, new_n7538,
    new_n7539, new_n7540, new_n7541, new_n7542, new_n7543, new_n7544,
    new_n7545, new_n7546, new_n7547, new_n7548, new_n7549, new_n7550,
    new_n7551, new_n7552, new_n7553, new_n7554, new_n7555, new_n7556,
    new_n7557, new_n7558, new_n7559, new_n7560, new_n7561, new_n7562,
    new_n7563, new_n7564, new_n7565, new_n7566, new_n7567, new_n7568,
    new_n7569, new_n7570, new_n7571, new_n7572, new_n7573, new_n7574,
    new_n7575, new_n7576, new_n7577, new_n7578, new_n7579, new_n7580,
    new_n7581, new_n7582, new_n7583, new_n7584, new_n7585, new_n7586,
    new_n7587, new_n7588, new_n7589, new_n7590, new_n7591, new_n7592,
    new_n7593, new_n7594, new_n7595, new_n7596, new_n7597, new_n7598,
    new_n7599, new_n7600, new_n7601, new_n7602, new_n7603, new_n7604,
    new_n7605, new_n7606, new_n7607, new_n7608, new_n7609, new_n7610,
    new_n7611, new_n7612, new_n7613, new_n7614, new_n7615, new_n7616,
    new_n7617, new_n7618, new_n7619, new_n7620, new_n7621, new_n7622,
    new_n7623, new_n7624, new_n7625, new_n7626, new_n7627, new_n7628,
    new_n7629, new_n7630, new_n7631, new_n7632, new_n7633, new_n7634,
    new_n7635, new_n7636, new_n7637, new_n7638, new_n7639, new_n7640,
    new_n7641, new_n7642, new_n7643, new_n7644, new_n7645, new_n7646,
    new_n7647, new_n7648, new_n7649, new_n7650, new_n7651, new_n7652,
    new_n7653, new_n7654, new_n7655, new_n7656, new_n7657, new_n7658,
    new_n7659, new_n7660, new_n7661, new_n7662, new_n7663, new_n7664,
    new_n7665, new_n7666, new_n7667, new_n7668, new_n7669, new_n7670,
    new_n7671, new_n7672, new_n7673, new_n7674, new_n7675, new_n7676,
    new_n7677, new_n7678, new_n7679, new_n7680, new_n7681, new_n7682,
    new_n7683, new_n7684, new_n7685, new_n7686, new_n7687, new_n7688,
    new_n7689, new_n7690, new_n7691, new_n7692, new_n7693, new_n7694,
    new_n7695, new_n7696, new_n7697, new_n7698, new_n7699, new_n7700,
    new_n7701, new_n7702, new_n7703, new_n7704, new_n7705, new_n7706,
    new_n7707, new_n7708, new_n7709, new_n7710, new_n7711, new_n7712,
    new_n7713, new_n7714, new_n7715, new_n7716, new_n7717, new_n7718,
    new_n7719, new_n7720, new_n7721, new_n7722, new_n7723, new_n7724,
    new_n7725, new_n7726, new_n7727, new_n7728, new_n7729, new_n7730,
    new_n7731, new_n7732, new_n7733, new_n7734, new_n7735, new_n7736,
    new_n7737, new_n7738, new_n7739, new_n7740, new_n7741, new_n7742,
    new_n7743, new_n7744, new_n7745, new_n7746, new_n7747, new_n7748,
    new_n7749, new_n7750, new_n7751, new_n7752, new_n7753, new_n7754,
    new_n7755, new_n7756, new_n7757, new_n7758, new_n7759, new_n7760,
    new_n7761, new_n7762, new_n7763, new_n7764, new_n7765, new_n7766,
    new_n7767, new_n7768, new_n7769, new_n7770, new_n7771, new_n7772,
    new_n7773, new_n7774, new_n7775, new_n7776, new_n7777, new_n7778,
    new_n7779, new_n7780, new_n7781, new_n7782, new_n7783, new_n7784,
    new_n7785, new_n7786, new_n7787, new_n7788, new_n7789, new_n7790,
    new_n7791, new_n7792, new_n7793, new_n7794, new_n7795, new_n7796,
    new_n7797, new_n7798, new_n7799, new_n7800, new_n7801, new_n7802,
    new_n7803, new_n7804, new_n7805, new_n7806, new_n7807, new_n7808,
    new_n7809, new_n7810, new_n7811, new_n7812, new_n7813, new_n7814,
    new_n7815, new_n7816, new_n7817, new_n7819, new_n7820, new_n7821,
    new_n7822, new_n7823, new_n7824, new_n7825, new_n7826, new_n7827,
    new_n7828, new_n7829, new_n7830, new_n7831, new_n7832, new_n7833,
    new_n7834, new_n7835, new_n7836, new_n7837, new_n7838, new_n7839,
    new_n7840, new_n7841, new_n7842, new_n7843, new_n7844, new_n7845,
    new_n7846, new_n7847, new_n7848, new_n7849, new_n7850, new_n7851,
    new_n7852, new_n7853, new_n7854, new_n7855, new_n7856, new_n7857,
    new_n7858, new_n7859, new_n7860, new_n7861, new_n7862, new_n7863,
    new_n7864, new_n7865, new_n7866, new_n7867, new_n7868, new_n7869,
    new_n7870, new_n7871, new_n7872, new_n7873, new_n7874, new_n7875,
    new_n7876, new_n7877, new_n7878, new_n7879, new_n7880, new_n7881,
    new_n7882, new_n7883, new_n7884, new_n7885, new_n7886, new_n7887,
    new_n7888, new_n7889, new_n7890, new_n7891, new_n7892, new_n7893,
    new_n7894, new_n7895, new_n7896, new_n7897, new_n7898, new_n7899,
    new_n7900, new_n7901, new_n7902, new_n7903, new_n7904, new_n7905,
    new_n7906, new_n7907, new_n7908, new_n7909, new_n7910, new_n7911,
    new_n7912, new_n7913, new_n7914, new_n7915, new_n7916, new_n7917,
    new_n7918, new_n7919, new_n7920, new_n7921, new_n7922, new_n7923,
    new_n7924, new_n7925, new_n7926, new_n7927, new_n7928, new_n7929,
    new_n7930, new_n7931, new_n7932, new_n7933, new_n7934, new_n7935,
    new_n7936, new_n7937, new_n7938, new_n7939, new_n7940, new_n7941,
    new_n7942, new_n7943, new_n7944, new_n7945, new_n7946, new_n7947,
    new_n7948, new_n7949, new_n7950, new_n7951, new_n7952, new_n7953,
    new_n7954, new_n7955, new_n7956, new_n7957, new_n7958, new_n7959,
    new_n7960, new_n7961, new_n7962, new_n7963, new_n7964, new_n7965,
    new_n7966, new_n7967, new_n7968, new_n7969, new_n7970, new_n7971,
    new_n7972, new_n7973, new_n7974, new_n7975, new_n7976, new_n7977,
    new_n7978, new_n7979, new_n7980, new_n7981, new_n7982, new_n7983,
    new_n7984, new_n7985, new_n7986, new_n7987, new_n7988, new_n7989,
    new_n7990, new_n7991, new_n7992, new_n7993, new_n7994, new_n7995,
    new_n7996, new_n7997, new_n7998, new_n7999, new_n8000, new_n8001,
    new_n8002, new_n8003, new_n8004, new_n8005, new_n8006, new_n8007,
    new_n8008, new_n8009, new_n8010, new_n8011, new_n8012, new_n8013,
    new_n8014, new_n8015, new_n8016, new_n8017, new_n8018, new_n8019,
    new_n8020, new_n8021, new_n8022, new_n8023, new_n8024, new_n8025,
    new_n8026, new_n8027, new_n8028, new_n8029, new_n8030, new_n8031,
    new_n8032, new_n8033, new_n8034, new_n8035, new_n8036, new_n8037,
    new_n8038, new_n8039, new_n8040, new_n8041, new_n8042, new_n8043,
    new_n8044, new_n8045, new_n8046, new_n8047, new_n8048, new_n8049,
    new_n8050, new_n8051, new_n8052, new_n8053, new_n8054, new_n8055,
    new_n8056, new_n8057, new_n8058, new_n8059, new_n8060, new_n8061,
    new_n8062, new_n8063, new_n8064, new_n8065, new_n8066, new_n8067,
    new_n8068, new_n8069, new_n8070, new_n8071, new_n8072, new_n8073,
    new_n8074, new_n8075, new_n8076, new_n8077, new_n8078, new_n8079,
    new_n8080, new_n8081, new_n8082, new_n8083, new_n8084, new_n8085,
    new_n8086, new_n8087, new_n8088, new_n8089, new_n8090, new_n8091,
    new_n8092, new_n8093, new_n8094, new_n8095, new_n8096, new_n8097,
    new_n8098, new_n8099, new_n8100, new_n8101, new_n8102, new_n8103,
    new_n8104, new_n8105, new_n8106, new_n8107, new_n8108, new_n8109,
    new_n8110, new_n8111, new_n8112, new_n8113, new_n8115, new_n8116,
    new_n8117, new_n8118, new_n8119, new_n8120, new_n8121, new_n8122,
    new_n8123, new_n8124, new_n8125, new_n8126, new_n8127, new_n8128,
    new_n8129, new_n8130, new_n8131, new_n8132, new_n8133, new_n8134,
    new_n8135, new_n8136, new_n8137, new_n8138, new_n8139, new_n8140,
    new_n8141, new_n8142, new_n8143, new_n8144, new_n8145, new_n8146,
    new_n8147, new_n8148, new_n8149, new_n8150, new_n8151, new_n8152,
    new_n8153, new_n8154, new_n8155, new_n8156, new_n8157, new_n8158,
    new_n8159, new_n8160, new_n8161, new_n8162, new_n8163, new_n8164,
    new_n8165, new_n8166, new_n8167, new_n8168, new_n8169, new_n8170,
    new_n8171, new_n8172, new_n8173, new_n8174, new_n8175, new_n8176,
    new_n8177, new_n8178, new_n8179, new_n8180, new_n8181, new_n8182,
    new_n8183, new_n8184, new_n8185, new_n8186, new_n8187, new_n8188,
    new_n8189, new_n8190, new_n8191, new_n8192, new_n8193, new_n8194,
    new_n8195, new_n8196, new_n8197, new_n8198, new_n8199, new_n8200,
    new_n8201, new_n8202, new_n8203, new_n8204, new_n8205, new_n8206,
    new_n8207, new_n8208, new_n8209, new_n8210, new_n8211, new_n8212,
    new_n8213, new_n8214, new_n8215, new_n8216, new_n8217, new_n8218,
    new_n8219, new_n8220, new_n8221, new_n8222, new_n8223, new_n8224,
    new_n8225, new_n8226, new_n8227, new_n8228, new_n8229, new_n8230,
    new_n8231, new_n8232, new_n8233, new_n8234, new_n8235, new_n8236,
    new_n8237, new_n8238, new_n8239, new_n8240, new_n8241, new_n8242,
    new_n8243, new_n8244, new_n8245, new_n8246, new_n8247, new_n8248,
    new_n8249, new_n8250, new_n8251, new_n8252, new_n8253, new_n8254,
    new_n8255, new_n8256, new_n8257, new_n8258, new_n8259, new_n8260,
    new_n8261, new_n8262, new_n8263, new_n8264, new_n8265, new_n8266,
    new_n8267, new_n8268, new_n8269, new_n8270, new_n8271, new_n8272,
    new_n8273, new_n8274, new_n8275, new_n8276, new_n8277, new_n8278,
    new_n8279, new_n8280, new_n8281, new_n8282, new_n8283, new_n8284,
    new_n8285, new_n8286, new_n8287, new_n8288, new_n8289, new_n8290,
    new_n8291, new_n8292, new_n8293, new_n8294, new_n8295, new_n8296,
    new_n8297, new_n8298, new_n8299, new_n8300, new_n8301, new_n8302,
    new_n8303, new_n8304, new_n8305, new_n8306, new_n8307, new_n8308,
    new_n8309, new_n8310, new_n8311, new_n8312, new_n8313, new_n8314,
    new_n8315, new_n8316, new_n8317, new_n8318, new_n8319, new_n8320,
    new_n8321, new_n8322, new_n8323, new_n8324, new_n8325, new_n8326,
    new_n8327, new_n8328, new_n8329, new_n8330, new_n8331, new_n8332,
    new_n8333, new_n8334, new_n8335, new_n8336, new_n8337, new_n8338,
    new_n8339, new_n8340, new_n8341, new_n8342, new_n8343, new_n8344,
    new_n8345, new_n8346, new_n8347, new_n8348, new_n8349, new_n8350,
    new_n8351, new_n8352, new_n8353, new_n8354, new_n8355, new_n8356,
    new_n8357, new_n8358, new_n8359, new_n8360, new_n8361, new_n8362,
    new_n8363, new_n8364, new_n8365, new_n8366, new_n8367, new_n8368,
    new_n8369, new_n8370, new_n8371, new_n8372, new_n8373, new_n8374,
    new_n8375, new_n8376, new_n8377, new_n8378, new_n8379, new_n8380,
    new_n8381, new_n8382, new_n8383, new_n8384, new_n8385, new_n8386,
    new_n8387, new_n8388, new_n8389, new_n8390, new_n8391, new_n8392,
    new_n8393, new_n8394, new_n8395, new_n8396, new_n8397, new_n8398,
    new_n8399, new_n8400, new_n8401, new_n8402, new_n8403, new_n8404,
    new_n8405, new_n8406, new_n8407, new_n8408, new_n8409, new_n8410,
    new_n8411, new_n8412, new_n8413, new_n8414, new_n8415, new_n8416,
    new_n8417, new_n8418, new_n8419, new_n8420, new_n8421, new_n8422,
    new_n8423, new_n8424, new_n8425, new_n8427, new_n8428, new_n8429,
    new_n8430, new_n8431, new_n8432, new_n8433, new_n8434, new_n8435,
    new_n8436, new_n8437, new_n8438, new_n8439, new_n8440, new_n8441,
    new_n8442, new_n8443, new_n8444, new_n8445, new_n8446, new_n8447,
    new_n8448, new_n8449, new_n8450, new_n8451, new_n8452, new_n8453,
    new_n8454, new_n8455, new_n8456, new_n8457, new_n8458, new_n8459,
    new_n8460, new_n8461, new_n8462, new_n8463, new_n8464, new_n8465,
    new_n8466, new_n8467, new_n8468, new_n8469, new_n8470, new_n8471,
    new_n8472, new_n8473, new_n8474, new_n8475, new_n8476, new_n8477,
    new_n8478, new_n8479, new_n8480, new_n8481, new_n8482, new_n8483,
    new_n8484, new_n8485, new_n8486, new_n8487, new_n8488, new_n8489,
    new_n8490, new_n8491, new_n8492, new_n8493, new_n8494, new_n8495,
    new_n8496, new_n8497, new_n8498, new_n8499, new_n8500, new_n8501,
    new_n8502, new_n8503, new_n8504, new_n8505, new_n8506, new_n8507,
    new_n8508, new_n8509, new_n8510, new_n8511, new_n8512, new_n8513,
    new_n8514, new_n8515, new_n8516, new_n8517, new_n8518, new_n8519,
    new_n8520, new_n8521, new_n8522, new_n8523, new_n8524, new_n8525,
    new_n8526, new_n8527, new_n8528, new_n8529, new_n8530, new_n8531,
    new_n8532, new_n8533, new_n8534, new_n8535, new_n8536, new_n8537,
    new_n8538, new_n8539, new_n8540, new_n8541, new_n8542, new_n8543,
    new_n8544, new_n8545, new_n8546, new_n8547, new_n8548, new_n8549,
    new_n8550, new_n8551, new_n8552, new_n8553, new_n8554, new_n8555,
    new_n8556, new_n8557, new_n8558, new_n8559, new_n8560, new_n8561,
    new_n8562, new_n8563, new_n8564, new_n8565, new_n8566, new_n8567,
    new_n8568, new_n8569, new_n8570, new_n8571, new_n8572, new_n8573,
    new_n8574, new_n8575, new_n8576, new_n8577, new_n8578, new_n8579,
    new_n8580, new_n8581, new_n8582, new_n8583, new_n8584, new_n8585,
    new_n8586, new_n8587, new_n8588, new_n8589, new_n8590, new_n8591,
    new_n8592, new_n8593, new_n8594, new_n8595, new_n8596, new_n8597,
    new_n8598, new_n8599, new_n8600, new_n8601, new_n8602, new_n8603,
    new_n8604, new_n8605, new_n8606, new_n8607, new_n8608, new_n8609,
    new_n8610, new_n8611, new_n8612, new_n8613, new_n8614, new_n8615,
    new_n8616, new_n8617, new_n8618, new_n8619, new_n8620, new_n8621,
    new_n8622, new_n8623, new_n8624, new_n8625, new_n8626, new_n8627,
    new_n8628, new_n8629, new_n8630, new_n8631, new_n8632, new_n8633,
    new_n8634, new_n8635, new_n8636, new_n8637, new_n8638, new_n8639,
    new_n8640, new_n8641, new_n8642, new_n8643, new_n8644, new_n8645,
    new_n8646, new_n8647, new_n8648, new_n8649, new_n8650, new_n8651,
    new_n8652, new_n8653, new_n8654, new_n8655, new_n8656, new_n8657,
    new_n8658, new_n8659, new_n8660, new_n8661, new_n8662, new_n8663,
    new_n8664, new_n8665, new_n8666, new_n8667, new_n8668, new_n8669,
    new_n8670, new_n8671, new_n8672, new_n8673, new_n8674, new_n8675,
    new_n8676, new_n8677, new_n8678, new_n8679, new_n8680, new_n8681,
    new_n8682, new_n8683, new_n8684, new_n8685, new_n8686, new_n8687,
    new_n8688, new_n8689, new_n8690, new_n8691, new_n8692, new_n8693,
    new_n8694, new_n8695, new_n8696, new_n8697, new_n8698, new_n8699,
    new_n8700, new_n8701, new_n8702, new_n8703, new_n8704, new_n8705,
    new_n8706, new_n8707, new_n8708, new_n8709, new_n8710, new_n8711,
    new_n8712, new_n8713, new_n8714, new_n8715, new_n8716, new_n8717,
    new_n8718, new_n8719, new_n8720, new_n8721, new_n8722, new_n8723,
    new_n8724, new_n8725, new_n8726, new_n8727, new_n8728, new_n8729,
    new_n8730, new_n8731, new_n8733, new_n8734, new_n8735, new_n8736,
    new_n8737, new_n8738, new_n8739, new_n8740, new_n8741, new_n8742,
    new_n8743, new_n8744, new_n8745, new_n8746, new_n8747, new_n8748,
    new_n8749, new_n8750, new_n8751, new_n8752, new_n8753, new_n8754,
    new_n8755, new_n8756, new_n8757, new_n8758, new_n8759, new_n8760,
    new_n8761, new_n8762, new_n8763, new_n8764, new_n8765, new_n8766,
    new_n8767, new_n8768, new_n8769, new_n8770, new_n8771, new_n8772,
    new_n8773, new_n8774, new_n8775, new_n8776, new_n8777, new_n8778,
    new_n8779, new_n8780, new_n8781, new_n8782, new_n8783, new_n8784,
    new_n8785, new_n8786, new_n8787, new_n8788, new_n8789, new_n8790,
    new_n8791, new_n8792, new_n8793, new_n8794, new_n8795, new_n8796,
    new_n8797, new_n8798, new_n8799, new_n8800, new_n8801, new_n8802,
    new_n8803, new_n8804, new_n8805, new_n8806, new_n8807, new_n8808,
    new_n8809, new_n8810, new_n8811, new_n8812, new_n8813, new_n8814,
    new_n8815, new_n8816, new_n8817, new_n8818, new_n8819, new_n8820,
    new_n8821, new_n8822, new_n8823, new_n8824, new_n8825, new_n8826,
    new_n8827, new_n8828, new_n8829, new_n8830, new_n8831, new_n8832,
    new_n8833, new_n8834, new_n8835, new_n8836, new_n8837, new_n8838,
    new_n8839, new_n8840, new_n8841, new_n8842, new_n8843, new_n8844,
    new_n8845, new_n8846, new_n8847, new_n8848, new_n8849, new_n8850,
    new_n8851, new_n8852, new_n8853, new_n8854, new_n8855, new_n8856,
    new_n8857, new_n8858, new_n8859, new_n8860, new_n8861, new_n8862,
    new_n8863, new_n8864, new_n8865, new_n8866, new_n8867, new_n8868,
    new_n8869, new_n8870, new_n8871, new_n8872, new_n8873, new_n8874,
    new_n8875, new_n8876, new_n8877, new_n8878, new_n8879, new_n8880,
    new_n8881, new_n8882, new_n8883, new_n8884, new_n8885, new_n8886,
    new_n8887, new_n8888, new_n8889, new_n8890, new_n8891, new_n8892,
    new_n8893, new_n8894, new_n8895, new_n8896, new_n8897, new_n8898,
    new_n8899, new_n8900, new_n8901, new_n8902, new_n8903, new_n8904,
    new_n8905, new_n8906, new_n8907, new_n8908, new_n8909, new_n8910,
    new_n8911, new_n8912, new_n8913, new_n8914, new_n8915, new_n8916,
    new_n8917, new_n8918, new_n8919, new_n8920, new_n8921, new_n8922,
    new_n8923, new_n8924, new_n8925, new_n8926, new_n8927, new_n8928,
    new_n8929, new_n8930, new_n8931, new_n8932, new_n8933, new_n8934,
    new_n8935, new_n8936, new_n8937, new_n8938, new_n8939, new_n8940,
    new_n8941, new_n8942, new_n8943, new_n8944, new_n8945, new_n8946,
    new_n8947, new_n8948, new_n8949, new_n8950, new_n8951, new_n8952,
    new_n8953, new_n8954, new_n8955, new_n8956, new_n8957, new_n8958,
    new_n8959, new_n8960, new_n8961, new_n8962, new_n8963, new_n8964,
    new_n8965, new_n8966, new_n8967, new_n8968, new_n8969, new_n8970,
    new_n8971, new_n8972, new_n8973, new_n8974, new_n8975, new_n8976,
    new_n8977, new_n8978, new_n8979, new_n8980, new_n8981, new_n8982,
    new_n8983, new_n8984, new_n8985, new_n8986, new_n8987, new_n8988,
    new_n8989, new_n8990, new_n8991, new_n8992, new_n8993, new_n8994,
    new_n8995, new_n8996, new_n8997, new_n8998, new_n8999, new_n9000,
    new_n9001, new_n9002, new_n9003, new_n9004, new_n9005, new_n9006,
    new_n9007, new_n9008, new_n9009, new_n9010, new_n9011, new_n9012,
    new_n9013, new_n9014, new_n9015, new_n9016, new_n9017, new_n9018,
    new_n9019, new_n9020, new_n9021, new_n9022, new_n9023, new_n9024,
    new_n9025, new_n9026, new_n9027, new_n9028, new_n9029, new_n9030,
    new_n9031, new_n9032, new_n9033, new_n9034, new_n9035, new_n9036,
    new_n9037, new_n9038, new_n9039, new_n9040, new_n9041, new_n9042,
    new_n9043, new_n9044, new_n9045, new_n9046, new_n9047, new_n9048,
    new_n9049, new_n9050, new_n9051, new_n9052, new_n9053, new_n9054,
    new_n9055, new_n9057, new_n9058, new_n9059, new_n9060, new_n9061,
    new_n9062, new_n9063, new_n9064, new_n9065, new_n9066, new_n9067,
    new_n9068, new_n9069, new_n9070, new_n9071, new_n9072, new_n9073,
    new_n9074, new_n9075, new_n9076, new_n9077, new_n9078, new_n9079,
    new_n9080, new_n9081, new_n9082, new_n9083, new_n9084, new_n9085,
    new_n9086, new_n9087, new_n9088, new_n9089, new_n9090, new_n9091,
    new_n9092, new_n9093, new_n9094, new_n9095, new_n9096, new_n9097,
    new_n9098, new_n9099, new_n9100, new_n9101, new_n9102, new_n9103,
    new_n9104, new_n9105, new_n9106, new_n9107, new_n9108, new_n9109,
    new_n9110, new_n9111, new_n9112, new_n9113, new_n9114, new_n9115,
    new_n9116, new_n9117, new_n9118, new_n9119, new_n9120, new_n9121,
    new_n9122, new_n9123, new_n9124, new_n9125, new_n9126, new_n9127,
    new_n9128, new_n9129, new_n9130, new_n9131, new_n9132, new_n9133,
    new_n9134, new_n9135, new_n9136, new_n9137, new_n9138, new_n9139,
    new_n9140, new_n9141, new_n9142, new_n9143, new_n9144, new_n9145,
    new_n9146, new_n9147, new_n9148, new_n9149, new_n9150, new_n9151,
    new_n9152, new_n9153, new_n9154, new_n9155, new_n9156, new_n9157,
    new_n9158, new_n9159, new_n9160, new_n9161, new_n9162, new_n9163,
    new_n9164, new_n9165, new_n9166, new_n9167, new_n9168, new_n9169,
    new_n9170, new_n9171, new_n9172, new_n9173, new_n9174, new_n9175,
    new_n9176, new_n9177, new_n9178, new_n9179, new_n9180, new_n9181,
    new_n9182, new_n9183, new_n9184, new_n9185, new_n9186, new_n9187,
    new_n9188, new_n9189, new_n9190, new_n9191, new_n9192, new_n9193,
    new_n9194, new_n9195, new_n9196, new_n9197, new_n9198, new_n9199,
    new_n9200, new_n9201, new_n9202, new_n9203, new_n9204, new_n9205,
    new_n9206, new_n9207, new_n9208, new_n9209, new_n9210, new_n9211,
    new_n9212, new_n9213, new_n9214, new_n9215, new_n9216, new_n9217,
    new_n9218, new_n9219, new_n9220, new_n9221, new_n9222, new_n9223,
    new_n9224, new_n9225, new_n9226, new_n9227, new_n9228, new_n9229,
    new_n9230, new_n9231, new_n9232, new_n9233, new_n9234, new_n9235,
    new_n9236, new_n9237, new_n9238, new_n9239, new_n9240, new_n9241,
    new_n9242, new_n9243, new_n9244, new_n9245, new_n9246, new_n9247,
    new_n9248, new_n9249, new_n9250, new_n9251, new_n9252, new_n9253,
    new_n9254, new_n9255, new_n9256, new_n9257, new_n9258, new_n9259,
    new_n9260, new_n9261, new_n9262, new_n9263, new_n9264, new_n9265,
    new_n9266, new_n9267, new_n9268, new_n9269, new_n9270, new_n9271,
    new_n9272, new_n9273, new_n9274, new_n9275, new_n9276, new_n9277,
    new_n9278, new_n9279, new_n9280, new_n9281, new_n9282, new_n9283,
    new_n9284, new_n9285, new_n9286, new_n9287, new_n9288, new_n9289,
    new_n9290, new_n9291, new_n9292, new_n9293, new_n9294, new_n9295,
    new_n9296, new_n9297, new_n9298, new_n9299, new_n9300, new_n9301,
    new_n9302, new_n9303, new_n9304, new_n9305, new_n9306, new_n9307,
    new_n9308, new_n9309, new_n9310, new_n9311, new_n9312, new_n9313,
    new_n9314, new_n9315, new_n9316, new_n9317, new_n9318, new_n9319,
    new_n9320, new_n9321, new_n9322, new_n9323, new_n9324, new_n9325,
    new_n9326, new_n9327, new_n9328, new_n9329, new_n9330, new_n9331,
    new_n9332, new_n9333, new_n9334, new_n9335, new_n9336, new_n9337,
    new_n9338, new_n9339, new_n9340, new_n9341, new_n9342, new_n9343,
    new_n9344, new_n9345, new_n9346, new_n9347, new_n9348, new_n9349,
    new_n9350, new_n9351, new_n9352, new_n9353, new_n9354, new_n9355,
    new_n9356, new_n9357, new_n9358, new_n9359, new_n9360, new_n9361,
    new_n9362, new_n9363, new_n9364, new_n9365, new_n9366, new_n9367,
    new_n9368, new_n9369, new_n9370, new_n9371, new_n9372, new_n9373,
    new_n9374, new_n9375, new_n9376, new_n9377, new_n9378, new_n9379,
    new_n9381, new_n9382, new_n9383, new_n9384, new_n9385, new_n9386,
    new_n9387, new_n9388, new_n9389, new_n9390, new_n9391, new_n9392,
    new_n9393, new_n9394, new_n9395, new_n9396, new_n9397, new_n9398,
    new_n9399, new_n9400, new_n9401, new_n9402, new_n9403, new_n9404,
    new_n9405, new_n9406, new_n9407, new_n9408, new_n9409, new_n9410,
    new_n9411, new_n9412, new_n9413, new_n9414, new_n9415, new_n9416,
    new_n9417, new_n9418, new_n9419, new_n9420, new_n9421, new_n9422,
    new_n9423, new_n9424, new_n9425, new_n9426, new_n9427, new_n9428,
    new_n9429, new_n9430, new_n9431, new_n9432, new_n9433, new_n9434,
    new_n9435, new_n9436, new_n9437, new_n9438, new_n9439, new_n9440,
    new_n9441, new_n9442, new_n9443, new_n9444, new_n9445, new_n9446,
    new_n9447, new_n9448, new_n9449, new_n9450, new_n9451, new_n9452,
    new_n9453, new_n9454, new_n9455, new_n9456, new_n9457, new_n9458,
    new_n9459, new_n9460, new_n9461, new_n9462, new_n9463, new_n9464,
    new_n9465, new_n9466, new_n9467, new_n9468, new_n9469, new_n9470,
    new_n9471, new_n9472, new_n9473, new_n9474, new_n9475, new_n9476,
    new_n9477, new_n9478, new_n9479, new_n9480, new_n9481, new_n9482,
    new_n9483, new_n9484, new_n9485, new_n9486, new_n9487, new_n9488,
    new_n9489, new_n9490, new_n9491, new_n9492, new_n9493, new_n9494,
    new_n9495, new_n9496, new_n9497, new_n9498, new_n9499, new_n9500,
    new_n9501, new_n9502, new_n9503, new_n9504, new_n9505, new_n9506,
    new_n9507, new_n9508, new_n9509, new_n9510, new_n9511, new_n9512,
    new_n9513, new_n9514, new_n9515, new_n9516, new_n9517, new_n9518,
    new_n9519, new_n9520, new_n9521, new_n9522, new_n9523, new_n9524,
    new_n9525, new_n9526, new_n9527, new_n9528, new_n9529, new_n9530,
    new_n9531, new_n9532, new_n9533, new_n9534, new_n9535, new_n9536,
    new_n9537, new_n9538, new_n9539, new_n9540, new_n9541, new_n9542,
    new_n9543, new_n9544, new_n9545, new_n9546, new_n9547, new_n9548,
    new_n9549, new_n9550, new_n9551, new_n9552, new_n9553, new_n9554,
    new_n9555, new_n9556, new_n9557, new_n9558, new_n9559, new_n9560,
    new_n9561, new_n9562, new_n9563, new_n9564, new_n9565, new_n9566,
    new_n9567, new_n9568, new_n9569, new_n9570, new_n9571, new_n9572,
    new_n9573, new_n9574, new_n9575, new_n9576, new_n9577, new_n9578,
    new_n9579, new_n9580, new_n9581, new_n9582, new_n9583, new_n9584,
    new_n9585, new_n9586, new_n9587, new_n9588, new_n9589, new_n9590,
    new_n9591, new_n9592, new_n9593, new_n9594, new_n9595, new_n9596,
    new_n9597, new_n9598, new_n9599, new_n9600, new_n9601, new_n9602,
    new_n9603, new_n9604, new_n9605, new_n9606, new_n9607, new_n9608,
    new_n9609, new_n9610, new_n9611, new_n9612, new_n9613, new_n9614,
    new_n9615, new_n9616, new_n9617, new_n9618, new_n9619, new_n9620,
    new_n9621, new_n9622, new_n9623, new_n9624, new_n9625, new_n9626,
    new_n9627, new_n9628, new_n9629, new_n9630, new_n9631, new_n9632,
    new_n9633, new_n9634, new_n9635, new_n9636, new_n9637, new_n9638,
    new_n9639, new_n9640, new_n9641, new_n9642, new_n9643, new_n9644,
    new_n9645, new_n9646, new_n9647, new_n9648, new_n9649, new_n9650,
    new_n9651, new_n9652, new_n9653, new_n9654, new_n9655, new_n9656,
    new_n9657, new_n9658, new_n9659, new_n9660, new_n9661, new_n9662,
    new_n9663, new_n9664, new_n9665, new_n9666, new_n9667, new_n9668,
    new_n9669, new_n9670, new_n9671, new_n9672, new_n9673, new_n9674,
    new_n9675, new_n9676, new_n9677, new_n9678, new_n9679, new_n9680,
    new_n9681, new_n9682, new_n9683, new_n9684, new_n9685, new_n9686,
    new_n9687, new_n9688, new_n9689, new_n9690, new_n9691, new_n9692,
    new_n9693, new_n9694, new_n9695, new_n9696, new_n9697, new_n9698,
    new_n9699, new_n9700, new_n9701, new_n9702, new_n9703, new_n9704,
    new_n9705, new_n9706, new_n9707, new_n9708, new_n9709, new_n9710,
    new_n9711, new_n9712, new_n9713, new_n9714, new_n9715, new_n9716,
    new_n9717, new_n9719, new_n9720, new_n9721, new_n9722, new_n9723,
    new_n9724, new_n9725, new_n9726, new_n9727, new_n9728, new_n9729,
    new_n9730, new_n9731, new_n9732, new_n9733, new_n9734, new_n9735,
    new_n9736, new_n9737, new_n9738, new_n9739, new_n9740, new_n9741,
    new_n9742, new_n9743, new_n9744, new_n9745, new_n9746, new_n9747,
    new_n9748, new_n9749, new_n9750, new_n9751, new_n9752, new_n9753,
    new_n9754, new_n9755, new_n9756, new_n9757, new_n9758, new_n9759,
    new_n9760, new_n9761, new_n9762, new_n9763, new_n9764, new_n9765,
    new_n9766, new_n9767, new_n9768, new_n9769, new_n9770, new_n9771,
    new_n9772, new_n9773, new_n9774, new_n9775, new_n9776, new_n9777,
    new_n9778, new_n9779, new_n9780, new_n9781, new_n9782, new_n9783,
    new_n9784, new_n9785, new_n9786, new_n9787, new_n9788, new_n9789,
    new_n9790, new_n9791, new_n9792, new_n9793, new_n9794, new_n9795,
    new_n9796, new_n9797, new_n9798, new_n9799, new_n9800, new_n9801,
    new_n9802, new_n9803, new_n9804, new_n9805, new_n9806, new_n9807,
    new_n9808, new_n9809, new_n9810, new_n9811, new_n9812, new_n9813,
    new_n9814, new_n9815, new_n9816, new_n9817, new_n9818, new_n9819,
    new_n9820, new_n9821, new_n9822, new_n9823, new_n9824, new_n9825,
    new_n9826, new_n9827, new_n9828, new_n9829, new_n9830, new_n9831,
    new_n9832, new_n9833, new_n9834, new_n9835, new_n9836, new_n9837,
    new_n9838, new_n9839, new_n9840, new_n9841, new_n9842, new_n9843,
    new_n9844, new_n9845, new_n9846, new_n9847, new_n9848, new_n9849,
    new_n9850, new_n9851, new_n9852, new_n9853, new_n9854, new_n9855,
    new_n9856, new_n9857, new_n9858, new_n9859, new_n9860, new_n9861,
    new_n9862, new_n9863, new_n9864, new_n9865, new_n9866, new_n9867,
    new_n9868, new_n9869, new_n9870, new_n9871, new_n9872, new_n9873,
    new_n9874, new_n9875, new_n9876, new_n9877, new_n9878, new_n9879,
    new_n9880, new_n9881, new_n9882, new_n9883, new_n9884, new_n9885,
    new_n9886, new_n9887, new_n9888, new_n9889, new_n9890, new_n9891,
    new_n9892, new_n9893, new_n9894, new_n9895, new_n9896, new_n9897,
    new_n9898, new_n9899, new_n9900, new_n9901, new_n9902, new_n9903,
    new_n9904, new_n9905, new_n9906, new_n9907, new_n9908, new_n9909,
    new_n9910, new_n9911, new_n9912, new_n9913, new_n9914, new_n9915,
    new_n9916, new_n9917, new_n9918, new_n9919, new_n9920, new_n9921,
    new_n9922, new_n9923, new_n9924, new_n9925, new_n9926, new_n9927,
    new_n9928, new_n9929, new_n9930, new_n9931, new_n9932, new_n9933,
    new_n9934, new_n9935, new_n9936, new_n9937, new_n9938, new_n9939,
    new_n9940, new_n9941, new_n9942, new_n9943, new_n9944, new_n9945,
    new_n9946, new_n9947, new_n9948, new_n9949, new_n9950, new_n9951,
    new_n9952, new_n9953, new_n9954, new_n9955, new_n9956, new_n9957,
    new_n9958, new_n9959, new_n9960, new_n9961, new_n9962, new_n9963,
    new_n9964, new_n9965, new_n9966, new_n9967, new_n9968, new_n9969,
    new_n9970, new_n9971, new_n9972, new_n9973, new_n9974, new_n9975,
    new_n9976, new_n9977, new_n9978, new_n9979, new_n9980, new_n9981,
    new_n9982, new_n9983, new_n9984, new_n9985, new_n9986, new_n9987,
    new_n9988, new_n9989, new_n9990, new_n9991, new_n9992, new_n9993,
    new_n9994, new_n9995, new_n9996, new_n9997, new_n9998, new_n9999,
    new_n10000, new_n10001, new_n10002, new_n10003, new_n10004, new_n10005,
    new_n10006, new_n10007, new_n10008, new_n10009, new_n10010, new_n10011,
    new_n10012, new_n10013, new_n10014, new_n10015, new_n10016, new_n10017,
    new_n10018, new_n10019, new_n10020, new_n10021, new_n10022, new_n10023,
    new_n10024, new_n10025, new_n10026, new_n10027, new_n10028, new_n10029,
    new_n10030, new_n10031, new_n10032, new_n10033, new_n10034, new_n10035,
    new_n10036, new_n10037, new_n10038, new_n10039, new_n10040, new_n10041,
    new_n10042, new_n10043, new_n10044, new_n10045, new_n10046, new_n10047,
    new_n10049, new_n10050, new_n10051, new_n10052, new_n10053, new_n10054,
    new_n10055, new_n10056, new_n10057, new_n10058, new_n10059, new_n10060,
    new_n10061, new_n10062, new_n10063, new_n10064, new_n10065, new_n10066,
    new_n10067, new_n10068, new_n10069, new_n10070, new_n10071, new_n10072,
    new_n10073, new_n10074, new_n10075, new_n10076, new_n10077, new_n10078,
    new_n10079, new_n10080, new_n10081, new_n10082, new_n10083, new_n10084,
    new_n10085, new_n10086, new_n10087, new_n10088, new_n10089, new_n10090,
    new_n10091, new_n10092, new_n10093, new_n10094, new_n10095, new_n10096,
    new_n10097, new_n10098, new_n10099, new_n10100, new_n10101, new_n10102,
    new_n10103, new_n10104, new_n10105, new_n10106, new_n10107, new_n10108,
    new_n10109, new_n10110, new_n10111, new_n10112, new_n10113, new_n10114,
    new_n10115, new_n10116, new_n10117, new_n10118, new_n10119, new_n10120,
    new_n10121, new_n10122, new_n10123, new_n10124, new_n10125, new_n10126,
    new_n10127, new_n10128, new_n10129, new_n10130, new_n10131, new_n10132,
    new_n10133, new_n10134, new_n10135, new_n10136, new_n10137, new_n10138,
    new_n10139, new_n10140, new_n10141, new_n10142, new_n10143, new_n10144,
    new_n10145, new_n10146, new_n10147, new_n10148, new_n10149, new_n10150,
    new_n10151, new_n10152, new_n10153, new_n10154, new_n10155, new_n10156,
    new_n10157, new_n10158, new_n10159, new_n10160, new_n10161, new_n10162,
    new_n10163, new_n10164, new_n10165, new_n10166, new_n10167, new_n10168,
    new_n10169, new_n10170, new_n10171, new_n10172, new_n10173, new_n10174,
    new_n10175, new_n10176, new_n10177, new_n10178, new_n10179, new_n10180,
    new_n10181, new_n10182, new_n10183, new_n10184, new_n10185, new_n10186,
    new_n10187, new_n10188, new_n10189, new_n10190, new_n10191, new_n10192,
    new_n10193, new_n10194, new_n10195, new_n10196, new_n10197, new_n10198,
    new_n10199, new_n10200, new_n10201, new_n10202, new_n10203, new_n10204,
    new_n10205, new_n10206, new_n10207, new_n10208, new_n10209, new_n10210,
    new_n10211, new_n10212, new_n10213, new_n10214, new_n10215, new_n10216,
    new_n10217, new_n10218, new_n10219, new_n10220, new_n10221, new_n10222,
    new_n10223, new_n10224, new_n10225, new_n10226, new_n10227, new_n10228,
    new_n10229, new_n10230, new_n10231, new_n10232, new_n10233, new_n10234,
    new_n10235, new_n10236, new_n10237, new_n10238, new_n10239, new_n10240,
    new_n10241, new_n10242, new_n10243, new_n10244, new_n10245, new_n10246,
    new_n10247, new_n10248, new_n10249, new_n10250, new_n10251, new_n10252,
    new_n10253, new_n10254, new_n10255, new_n10256, new_n10257, new_n10258,
    new_n10259, new_n10260, new_n10261, new_n10262, new_n10263, new_n10264,
    new_n10265, new_n10266, new_n10267, new_n10268, new_n10269, new_n10270,
    new_n10271, new_n10272, new_n10273, new_n10274, new_n10275, new_n10276,
    new_n10277, new_n10278, new_n10279, new_n10280, new_n10281, new_n10282,
    new_n10283, new_n10284, new_n10285, new_n10286, new_n10287, new_n10288,
    new_n10289, new_n10290, new_n10291, new_n10292, new_n10293, new_n10294,
    new_n10295, new_n10296, new_n10297, new_n10298, new_n10299, new_n10300,
    new_n10301, new_n10302, new_n10303, new_n10304, new_n10305, new_n10306,
    new_n10307, new_n10308, new_n10309, new_n10310, new_n10311, new_n10312,
    new_n10313, new_n10314, new_n10315, new_n10316, new_n10317, new_n10318,
    new_n10319, new_n10320, new_n10321, new_n10322, new_n10323, new_n10324,
    new_n10325, new_n10326, new_n10327, new_n10328, new_n10329, new_n10330,
    new_n10331, new_n10332, new_n10333, new_n10334, new_n10335, new_n10336,
    new_n10337, new_n10338, new_n10339, new_n10340, new_n10341, new_n10342,
    new_n10343, new_n10344, new_n10345, new_n10346, new_n10347, new_n10348,
    new_n10349, new_n10350, new_n10351, new_n10352, new_n10353, new_n10354,
    new_n10355, new_n10356, new_n10357, new_n10358, new_n10359, new_n10360,
    new_n10361, new_n10362, new_n10363, new_n10364, new_n10365, new_n10366,
    new_n10367, new_n10368, new_n10369, new_n10370, new_n10371, new_n10372,
    new_n10373, new_n10374, new_n10375, new_n10376, new_n10377, new_n10378,
    new_n10379, new_n10380, new_n10381, new_n10382, new_n10383, new_n10384,
    new_n10385, new_n10386, new_n10387, new_n10388, new_n10389, new_n10390,
    new_n10391, new_n10392, new_n10393, new_n10394, new_n10395, new_n10397,
    new_n10398, new_n10399, new_n10400, new_n10401, new_n10402, new_n10403,
    new_n10404, new_n10405, new_n10406, new_n10407, new_n10408, new_n10409,
    new_n10410, new_n10411, new_n10412, new_n10413, new_n10414, new_n10415,
    new_n10416, new_n10417, new_n10418, new_n10419, new_n10420, new_n10421,
    new_n10422, new_n10423, new_n10424, new_n10425, new_n10426, new_n10427,
    new_n10428, new_n10429, new_n10430, new_n10431, new_n10432, new_n10433,
    new_n10434, new_n10435, new_n10436, new_n10437, new_n10438, new_n10439,
    new_n10440, new_n10441, new_n10442, new_n10443, new_n10444, new_n10445,
    new_n10446, new_n10447, new_n10448, new_n10449, new_n10450, new_n10451,
    new_n10452, new_n10453, new_n10454, new_n10455, new_n10456, new_n10457,
    new_n10458, new_n10459, new_n10460, new_n10461, new_n10462, new_n10463,
    new_n10464, new_n10465, new_n10466, new_n10467, new_n10468, new_n10469,
    new_n10470, new_n10471, new_n10472, new_n10473, new_n10474, new_n10475,
    new_n10476, new_n10477, new_n10478, new_n10479, new_n10480, new_n10481,
    new_n10482, new_n10483, new_n10484, new_n10485, new_n10486, new_n10487,
    new_n10488, new_n10489, new_n10490, new_n10491, new_n10492, new_n10493,
    new_n10494, new_n10495, new_n10496, new_n10497, new_n10498, new_n10499,
    new_n10500, new_n10501, new_n10502, new_n10503, new_n10504, new_n10505,
    new_n10506, new_n10507, new_n10508, new_n10509, new_n10510, new_n10511,
    new_n10512, new_n10513, new_n10514, new_n10515, new_n10516, new_n10517,
    new_n10518, new_n10519, new_n10520, new_n10521, new_n10522, new_n10523,
    new_n10524, new_n10525, new_n10526, new_n10527, new_n10528, new_n10529,
    new_n10530, new_n10531, new_n10532, new_n10533, new_n10534, new_n10535,
    new_n10536, new_n10537, new_n10538, new_n10539, new_n10540, new_n10541,
    new_n10542, new_n10543, new_n10544, new_n10545, new_n10546, new_n10547,
    new_n10548, new_n10549, new_n10550, new_n10551, new_n10552, new_n10553,
    new_n10554, new_n10555, new_n10556, new_n10557, new_n10558, new_n10559,
    new_n10560, new_n10561, new_n10562, new_n10563, new_n10564, new_n10565,
    new_n10566, new_n10567, new_n10568, new_n10569, new_n10570, new_n10571,
    new_n10572, new_n10573, new_n10574, new_n10575, new_n10576, new_n10577,
    new_n10578, new_n10579, new_n10580, new_n10581, new_n10582, new_n10583,
    new_n10584, new_n10585, new_n10586, new_n10587, new_n10588, new_n10589,
    new_n10590, new_n10591, new_n10592, new_n10593, new_n10594, new_n10595,
    new_n10596, new_n10597, new_n10598, new_n10599, new_n10600, new_n10601,
    new_n10602, new_n10603, new_n10604, new_n10605, new_n10606, new_n10607,
    new_n10608, new_n10609, new_n10610, new_n10611, new_n10612, new_n10613,
    new_n10614, new_n10615, new_n10616, new_n10617, new_n10618, new_n10619,
    new_n10620, new_n10621, new_n10622, new_n10623, new_n10624, new_n10625,
    new_n10626, new_n10627, new_n10628, new_n10629, new_n10630, new_n10631,
    new_n10632, new_n10633, new_n10634, new_n10635, new_n10636, new_n10637,
    new_n10638, new_n10639, new_n10640, new_n10641, new_n10642, new_n10643,
    new_n10644, new_n10645, new_n10646, new_n10647, new_n10648, new_n10649,
    new_n10650, new_n10651, new_n10652, new_n10653, new_n10654, new_n10655,
    new_n10656, new_n10657, new_n10658, new_n10659, new_n10660, new_n10661,
    new_n10662, new_n10663, new_n10664, new_n10665, new_n10666, new_n10667,
    new_n10668, new_n10669, new_n10670, new_n10671, new_n10672, new_n10673,
    new_n10674, new_n10675, new_n10676, new_n10677, new_n10678, new_n10679,
    new_n10680, new_n10681, new_n10682, new_n10683, new_n10684, new_n10685,
    new_n10686, new_n10687, new_n10688, new_n10689, new_n10690, new_n10691,
    new_n10692, new_n10693, new_n10694, new_n10695, new_n10696, new_n10697,
    new_n10698, new_n10699, new_n10700, new_n10701, new_n10702, new_n10703,
    new_n10704, new_n10705, new_n10706, new_n10707, new_n10708, new_n10709,
    new_n10710, new_n10711, new_n10712, new_n10713, new_n10714, new_n10715,
    new_n10716, new_n10717, new_n10718, new_n10719, new_n10720, new_n10721,
    new_n10722, new_n10723, new_n10724, new_n10725, new_n10726, new_n10727,
    new_n10728, new_n10729, new_n10730, new_n10731, new_n10732, new_n10733,
    new_n10734, new_n10735, new_n10736, new_n10737, new_n10738, new_n10739,
    new_n10740, new_n10741, new_n10742, new_n10743, new_n10744, new_n10745,
    new_n10747, new_n10748, new_n10749, new_n10750, new_n10751, new_n10752,
    new_n10753, new_n10754, new_n10755, new_n10756, new_n10757, new_n10758,
    new_n10759, new_n10760, new_n10761, new_n10762, new_n10763, new_n10764,
    new_n10765, new_n10766, new_n10767, new_n10768, new_n10769, new_n10770,
    new_n10771, new_n10772, new_n10773, new_n10774, new_n10775, new_n10776,
    new_n10777, new_n10778, new_n10779, new_n10780, new_n10781, new_n10782,
    new_n10783, new_n10784, new_n10785, new_n10786, new_n10787, new_n10788,
    new_n10789, new_n10790, new_n10791, new_n10792, new_n10793, new_n10794,
    new_n10795, new_n10796, new_n10797, new_n10798, new_n10799, new_n10800,
    new_n10801, new_n10802, new_n10803, new_n10804, new_n10805, new_n10806,
    new_n10807, new_n10808, new_n10809, new_n10810, new_n10811, new_n10812,
    new_n10813, new_n10814, new_n10815, new_n10816, new_n10817, new_n10818,
    new_n10819, new_n10820, new_n10821, new_n10822, new_n10823, new_n10824,
    new_n10825, new_n10826, new_n10827, new_n10828, new_n10829, new_n10830,
    new_n10831, new_n10832, new_n10833, new_n10834, new_n10835, new_n10836,
    new_n10837, new_n10838, new_n10839, new_n10840, new_n10841, new_n10842,
    new_n10843, new_n10844, new_n10845, new_n10846, new_n10847, new_n10848,
    new_n10849, new_n10850, new_n10851, new_n10852, new_n10853, new_n10854,
    new_n10855, new_n10856, new_n10857, new_n10858, new_n10859, new_n10860,
    new_n10861, new_n10862, new_n10863, new_n10864, new_n10865, new_n10866,
    new_n10867, new_n10868, new_n10869, new_n10870, new_n10871, new_n10872,
    new_n10873, new_n10874, new_n10875, new_n10876, new_n10877, new_n10878,
    new_n10879, new_n10880, new_n10881, new_n10882, new_n10883, new_n10884,
    new_n10885, new_n10886, new_n10887, new_n10888, new_n10889, new_n10890,
    new_n10891, new_n10892, new_n10893, new_n10894, new_n10895, new_n10896,
    new_n10897, new_n10898, new_n10899, new_n10900, new_n10901, new_n10902,
    new_n10903, new_n10904, new_n10905, new_n10906, new_n10907, new_n10908,
    new_n10909, new_n10910, new_n10911, new_n10912, new_n10913, new_n10914,
    new_n10915, new_n10916, new_n10917, new_n10918, new_n10919, new_n10920,
    new_n10921, new_n10922, new_n10923, new_n10924, new_n10925, new_n10926,
    new_n10927, new_n10928, new_n10929, new_n10930, new_n10931, new_n10932,
    new_n10933, new_n10934, new_n10935, new_n10936, new_n10937, new_n10938,
    new_n10939, new_n10940, new_n10941, new_n10942, new_n10943, new_n10944,
    new_n10945, new_n10946, new_n10947, new_n10948, new_n10949, new_n10950,
    new_n10951, new_n10952, new_n10953, new_n10954, new_n10955, new_n10956,
    new_n10957, new_n10958, new_n10959, new_n10960, new_n10961, new_n10962,
    new_n10963, new_n10964, new_n10965, new_n10966, new_n10967, new_n10968,
    new_n10969, new_n10970, new_n10971, new_n10972, new_n10973, new_n10974,
    new_n10975, new_n10976, new_n10977, new_n10978, new_n10979, new_n10980,
    new_n10981, new_n10982, new_n10983, new_n10984, new_n10985, new_n10986,
    new_n10987, new_n10988, new_n10989, new_n10990, new_n10991, new_n10992,
    new_n10993, new_n10994, new_n10995, new_n10996, new_n10997, new_n10998,
    new_n10999, new_n11000, new_n11001, new_n11002, new_n11003, new_n11004,
    new_n11005, new_n11006, new_n11007, new_n11008, new_n11009, new_n11010,
    new_n11011, new_n11012, new_n11013, new_n11014, new_n11015, new_n11016,
    new_n11017, new_n11018, new_n11019, new_n11020, new_n11021, new_n11022,
    new_n11023, new_n11024, new_n11025, new_n11026, new_n11027, new_n11028,
    new_n11029, new_n11030, new_n11031, new_n11032, new_n11033, new_n11034,
    new_n11035, new_n11036, new_n11037, new_n11038, new_n11039, new_n11040,
    new_n11041, new_n11042, new_n11043, new_n11044, new_n11045, new_n11046,
    new_n11047, new_n11048, new_n11049, new_n11050, new_n11051, new_n11052,
    new_n11053, new_n11054, new_n11055, new_n11056, new_n11057, new_n11058,
    new_n11059, new_n11060, new_n11061, new_n11062, new_n11063, new_n11064,
    new_n11065, new_n11066, new_n11067, new_n11068, new_n11069, new_n11070,
    new_n11071, new_n11072, new_n11073, new_n11074, new_n11075, new_n11076,
    new_n11077, new_n11078, new_n11079, new_n11080, new_n11081, new_n11082,
    new_n11083, new_n11084, new_n11085, new_n11086, new_n11087, new_n11088,
    new_n11089, new_n11090, new_n11091, new_n11092, new_n11093, new_n11094,
    new_n11095, new_n11096, new_n11097, new_n11098, new_n11099, new_n11100,
    new_n11101, new_n11103, new_n11104, new_n11105, new_n11106, new_n11107,
    new_n11108, new_n11109, new_n11110, new_n11111, new_n11112, new_n11113,
    new_n11114, new_n11115, new_n11116, new_n11117, new_n11118, new_n11119,
    new_n11120, new_n11121, new_n11122, new_n11123, new_n11124, new_n11125,
    new_n11126, new_n11127, new_n11128, new_n11129, new_n11130, new_n11131,
    new_n11132, new_n11133, new_n11134, new_n11135, new_n11136, new_n11137,
    new_n11138, new_n11139, new_n11140, new_n11141, new_n11142, new_n11143,
    new_n11144, new_n11145, new_n11146, new_n11147, new_n11148, new_n11149,
    new_n11150, new_n11151, new_n11152, new_n11153, new_n11154, new_n11155,
    new_n11156, new_n11157, new_n11158, new_n11159, new_n11160, new_n11161,
    new_n11162, new_n11163, new_n11164, new_n11165, new_n11166, new_n11167,
    new_n11168, new_n11169, new_n11170, new_n11171, new_n11172, new_n11173,
    new_n11174, new_n11175, new_n11176, new_n11177, new_n11178, new_n11179,
    new_n11180, new_n11181, new_n11182, new_n11183, new_n11184, new_n11185,
    new_n11186, new_n11187, new_n11188, new_n11189, new_n11190, new_n11191,
    new_n11192, new_n11193, new_n11194, new_n11195, new_n11196, new_n11197,
    new_n11198, new_n11199, new_n11200, new_n11201, new_n11202, new_n11203,
    new_n11204, new_n11205, new_n11206, new_n11207, new_n11208, new_n11209,
    new_n11210, new_n11211, new_n11212, new_n11213, new_n11214, new_n11215,
    new_n11216, new_n11217, new_n11218, new_n11219, new_n11220, new_n11221,
    new_n11222, new_n11223, new_n11224, new_n11225, new_n11226, new_n11227,
    new_n11228, new_n11229, new_n11230, new_n11231, new_n11232, new_n11233,
    new_n11234, new_n11235, new_n11236, new_n11237, new_n11238, new_n11239,
    new_n11240, new_n11241, new_n11242, new_n11243, new_n11244, new_n11245,
    new_n11246, new_n11247, new_n11248, new_n11249, new_n11250, new_n11251,
    new_n11252, new_n11253, new_n11254, new_n11255, new_n11256, new_n11257,
    new_n11258, new_n11259, new_n11260, new_n11261, new_n11262, new_n11263,
    new_n11264, new_n11265, new_n11266, new_n11267, new_n11268, new_n11269,
    new_n11270, new_n11271, new_n11272, new_n11273, new_n11274, new_n11275,
    new_n11276, new_n11277, new_n11278, new_n11279, new_n11280, new_n11281,
    new_n11282, new_n11283, new_n11284, new_n11285, new_n11286, new_n11287,
    new_n11288, new_n11289, new_n11290, new_n11291, new_n11292, new_n11293,
    new_n11294, new_n11295, new_n11296, new_n11297, new_n11298, new_n11299,
    new_n11300, new_n11301, new_n11302, new_n11303, new_n11304, new_n11305,
    new_n11306, new_n11307, new_n11308, new_n11309, new_n11310, new_n11311,
    new_n11312, new_n11313, new_n11314, new_n11315, new_n11316, new_n11317,
    new_n11318, new_n11319, new_n11320, new_n11321, new_n11322, new_n11323,
    new_n11324, new_n11325, new_n11326, new_n11327, new_n11328, new_n11329,
    new_n11330, new_n11331, new_n11332, new_n11333, new_n11334, new_n11335,
    new_n11336, new_n11337, new_n11338, new_n11339, new_n11340, new_n11341,
    new_n11342, new_n11343, new_n11344, new_n11345, new_n11346, new_n11347,
    new_n11348, new_n11349, new_n11350, new_n11351, new_n11352, new_n11353,
    new_n11354, new_n11355, new_n11356, new_n11357, new_n11358, new_n11359,
    new_n11360, new_n11361, new_n11362, new_n11363, new_n11364, new_n11365,
    new_n11366, new_n11367, new_n11368, new_n11369, new_n11370, new_n11371,
    new_n11372, new_n11373, new_n11374, new_n11375, new_n11376, new_n11377,
    new_n11378, new_n11379, new_n11380, new_n11381, new_n11382, new_n11383,
    new_n11384, new_n11385, new_n11386, new_n11387, new_n11388, new_n11389,
    new_n11390, new_n11391, new_n11392, new_n11393, new_n11394, new_n11395,
    new_n11396, new_n11397, new_n11398, new_n11399, new_n11400, new_n11401,
    new_n11402, new_n11403, new_n11404, new_n11405, new_n11406, new_n11407,
    new_n11408, new_n11409, new_n11410, new_n11411, new_n11412, new_n11413,
    new_n11414, new_n11415, new_n11416, new_n11417, new_n11418, new_n11419,
    new_n11420, new_n11421, new_n11422, new_n11423, new_n11424, new_n11425,
    new_n11426, new_n11427, new_n11428, new_n11429, new_n11430, new_n11431,
    new_n11432, new_n11433, new_n11434, new_n11435, new_n11436, new_n11437,
    new_n11438, new_n11439, new_n11440, new_n11441, new_n11442, new_n11443,
    new_n11444, new_n11445, new_n11446, new_n11447, new_n11448, new_n11449,
    new_n11450, new_n11451, new_n11452, new_n11453, new_n11454, new_n11455,
    new_n11456, new_n11457, new_n11458, new_n11459, new_n11461, new_n11462,
    new_n11463, new_n11464, new_n11465, new_n11466, new_n11467, new_n11468,
    new_n11469, new_n11470, new_n11471, new_n11472, new_n11473, new_n11474,
    new_n11475, new_n11476, new_n11477, new_n11478, new_n11479, new_n11480,
    new_n11481, new_n11482, new_n11483, new_n11484, new_n11485, new_n11486,
    new_n11487, new_n11488, new_n11489, new_n11490, new_n11491, new_n11492,
    new_n11493, new_n11494, new_n11495, new_n11496, new_n11497, new_n11498,
    new_n11499, new_n11500, new_n11501, new_n11502, new_n11503, new_n11504,
    new_n11505, new_n11506, new_n11507, new_n11508, new_n11509, new_n11510,
    new_n11511, new_n11512, new_n11513, new_n11514, new_n11515, new_n11516,
    new_n11517, new_n11518, new_n11519, new_n11520, new_n11521, new_n11522,
    new_n11523, new_n11524, new_n11525, new_n11526, new_n11527, new_n11528,
    new_n11529, new_n11530, new_n11531, new_n11532, new_n11533, new_n11534,
    new_n11535, new_n11536, new_n11537, new_n11538, new_n11539, new_n11540,
    new_n11541, new_n11542, new_n11543, new_n11544, new_n11545, new_n11546,
    new_n11547, new_n11548, new_n11549, new_n11550, new_n11551, new_n11552,
    new_n11553, new_n11554, new_n11555, new_n11556, new_n11557, new_n11558,
    new_n11559, new_n11560, new_n11561, new_n11562, new_n11563, new_n11564,
    new_n11565, new_n11566, new_n11567, new_n11568, new_n11569, new_n11570,
    new_n11571, new_n11572, new_n11573, new_n11574, new_n11575, new_n11576,
    new_n11577, new_n11578, new_n11579, new_n11580, new_n11581, new_n11582,
    new_n11583, new_n11584, new_n11585, new_n11586, new_n11587, new_n11588,
    new_n11589, new_n11590, new_n11591, new_n11592, new_n11593, new_n11594,
    new_n11595, new_n11596, new_n11597, new_n11598, new_n11599, new_n11600,
    new_n11601, new_n11602, new_n11603, new_n11604, new_n11605, new_n11606,
    new_n11607, new_n11608, new_n11609, new_n11610, new_n11611, new_n11612,
    new_n11613, new_n11614, new_n11615, new_n11616, new_n11617, new_n11618,
    new_n11619, new_n11620, new_n11621, new_n11622, new_n11623, new_n11624,
    new_n11625, new_n11626, new_n11627, new_n11628, new_n11629, new_n11630,
    new_n11631, new_n11632, new_n11633, new_n11634, new_n11635, new_n11636,
    new_n11637, new_n11638, new_n11639, new_n11640, new_n11641, new_n11642,
    new_n11643, new_n11644, new_n11645, new_n11646, new_n11647, new_n11648,
    new_n11649, new_n11650, new_n11651, new_n11652, new_n11653, new_n11654,
    new_n11655, new_n11656, new_n11657, new_n11658, new_n11659, new_n11660,
    new_n11661, new_n11662, new_n11663, new_n11664, new_n11665, new_n11666,
    new_n11667, new_n11668, new_n11669, new_n11670, new_n11671, new_n11672,
    new_n11673, new_n11674, new_n11675, new_n11676, new_n11677, new_n11678,
    new_n11679, new_n11680, new_n11681, new_n11682, new_n11683, new_n11684,
    new_n11685, new_n11686, new_n11687, new_n11688, new_n11689, new_n11690,
    new_n11691, new_n11692, new_n11693, new_n11694, new_n11695, new_n11696,
    new_n11697, new_n11698, new_n11699, new_n11700, new_n11701, new_n11702,
    new_n11703, new_n11704, new_n11705, new_n11706, new_n11707, new_n11708,
    new_n11709, new_n11710, new_n11711, new_n11712, new_n11713, new_n11714,
    new_n11715, new_n11716, new_n11717, new_n11718, new_n11719, new_n11720,
    new_n11721, new_n11722, new_n11723, new_n11724, new_n11725, new_n11726,
    new_n11727, new_n11728, new_n11729, new_n11730, new_n11731, new_n11732,
    new_n11733, new_n11734, new_n11735, new_n11736, new_n11737, new_n11738,
    new_n11739, new_n11740, new_n11741, new_n11742, new_n11743, new_n11744,
    new_n11745, new_n11746, new_n11747, new_n11748, new_n11749, new_n11750,
    new_n11751, new_n11752, new_n11753, new_n11754, new_n11755, new_n11756,
    new_n11757, new_n11758, new_n11759, new_n11760, new_n11761, new_n11762,
    new_n11763, new_n11764, new_n11765, new_n11766, new_n11767, new_n11768,
    new_n11769, new_n11770, new_n11771, new_n11772, new_n11773, new_n11774,
    new_n11775, new_n11776, new_n11777, new_n11778, new_n11779, new_n11780,
    new_n11781, new_n11782, new_n11783, new_n11784, new_n11785, new_n11786,
    new_n11787, new_n11788, new_n11789, new_n11790, new_n11791, new_n11792,
    new_n11793, new_n11794, new_n11795, new_n11796, new_n11797, new_n11798,
    new_n11799, new_n11800, new_n11801, new_n11802, new_n11803, new_n11804,
    new_n11805, new_n11806, new_n11807, new_n11808, new_n11809, new_n11810,
    new_n11811, new_n11812, new_n11813, new_n11814, new_n11815, new_n11816,
    new_n11817, new_n11818, new_n11819, new_n11820, new_n11821, new_n11822,
    new_n11823, new_n11824, new_n11825, new_n11827, new_n11828, new_n11829,
    new_n11830, new_n11831, new_n11832, new_n11833, new_n11834, new_n11835,
    new_n11836, new_n11837, new_n11838, new_n11839, new_n11840, new_n11841,
    new_n11842, new_n11843, new_n11844, new_n11845, new_n11846, new_n11847,
    new_n11848, new_n11849, new_n11850, new_n11851, new_n11852, new_n11853,
    new_n11854, new_n11855, new_n11856, new_n11857, new_n11858, new_n11859,
    new_n11860, new_n11861, new_n11862, new_n11863, new_n11864, new_n11865,
    new_n11866, new_n11867, new_n11868, new_n11869, new_n11870, new_n11871,
    new_n11872, new_n11873, new_n11874, new_n11875, new_n11876, new_n11877,
    new_n11878, new_n11879, new_n11880, new_n11881, new_n11882, new_n11883,
    new_n11884, new_n11885, new_n11886, new_n11887, new_n11888, new_n11889,
    new_n11890, new_n11891, new_n11892, new_n11893, new_n11894, new_n11895,
    new_n11896, new_n11897, new_n11898, new_n11899, new_n11900, new_n11901,
    new_n11902, new_n11903, new_n11904, new_n11905, new_n11906, new_n11907,
    new_n11908, new_n11909, new_n11910, new_n11911, new_n11912, new_n11913,
    new_n11914, new_n11915, new_n11916, new_n11917, new_n11918, new_n11919,
    new_n11920, new_n11921, new_n11922, new_n11923, new_n11924, new_n11925,
    new_n11926, new_n11927, new_n11928, new_n11929, new_n11930, new_n11931,
    new_n11932, new_n11933, new_n11934, new_n11935, new_n11936, new_n11937,
    new_n11938, new_n11939, new_n11940, new_n11941, new_n11942, new_n11943,
    new_n11944, new_n11945, new_n11946, new_n11947, new_n11948, new_n11949,
    new_n11950, new_n11951, new_n11952, new_n11953, new_n11954, new_n11955,
    new_n11956, new_n11957, new_n11958, new_n11959, new_n11960, new_n11961,
    new_n11962, new_n11963, new_n11964, new_n11965, new_n11966, new_n11967,
    new_n11968, new_n11969, new_n11970, new_n11971, new_n11972, new_n11973,
    new_n11974, new_n11975, new_n11976, new_n11977, new_n11978, new_n11979,
    new_n11980, new_n11981, new_n11982, new_n11983, new_n11984, new_n11985,
    new_n11986, new_n11987, new_n11988, new_n11989, new_n11990, new_n11991,
    new_n11992, new_n11993, new_n11994, new_n11995, new_n11996, new_n11997,
    new_n11998, new_n11999, new_n12000, new_n12001, new_n12002, new_n12003,
    new_n12004, new_n12005, new_n12006, new_n12007, new_n12008, new_n12009,
    new_n12010, new_n12011, new_n12012, new_n12013, new_n12014, new_n12015,
    new_n12016, new_n12017, new_n12018, new_n12019, new_n12020, new_n12021,
    new_n12022, new_n12023, new_n12024, new_n12025, new_n12026, new_n12027,
    new_n12028, new_n12029, new_n12030, new_n12031, new_n12032, new_n12033,
    new_n12034, new_n12035, new_n12036, new_n12037, new_n12038, new_n12039,
    new_n12040, new_n12041, new_n12042, new_n12043, new_n12044, new_n12045,
    new_n12046, new_n12047, new_n12048, new_n12049, new_n12050, new_n12051,
    new_n12052, new_n12053, new_n12054, new_n12055, new_n12056, new_n12057,
    new_n12058, new_n12059, new_n12060, new_n12061, new_n12062, new_n12063,
    new_n12064, new_n12065, new_n12066, new_n12067, new_n12068, new_n12069,
    new_n12070, new_n12071, new_n12072, new_n12073, new_n12074, new_n12075,
    new_n12076, new_n12077, new_n12078, new_n12079, new_n12080, new_n12081,
    new_n12082, new_n12083, new_n12084, new_n12085, new_n12086, new_n12087,
    new_n12088, new_n12089, new_n12090, new_n12091, new_n12092, new_n12093,
    new_n12094, new_n12095, new_n12096, new_n12097, new_n12098, new_n12099,
    new_n12100, new_n12101, new_n12102, new_n12103, new_n12104, new_n12105,
    new_n12106, new_n12107, new_n12108, new_n12109, new_n12110, new_n12111,
    new_n12112, new_n12113, new_n12114, new_n12115, new_n12116, new_n12117,
    new_n12118, new_n12119, new_n12120, new_n12121, new_n12122, new_n12123,
    new_n12124, new_n12125, new_n12126, new_n12127, new_n12128, new_n12129,
    new_n12130, new_n12131, new_n12132, new_n12133, new_n12134, new_n12135,
    new_n12136, new_n12137, new_n12138, new_n12139, new_n12140, new_n12141,
    new_n12142, new_n12143, new_n12144, new_n12145, new_n12146, new_n12147,
    new_n12148, new_n12149, new_n12150, new_n12151, new_n12152, new_n12153,
    new_n12154, new_n12155, new_n12156, new_n12157, new_n12158, new_n12159,
    new_n12160, new_n12161, new_n12162, new_n12163, new_n12164, new_n12165,
    new_n12166, new_n12167, new_n12168, new_n12169, new_n12170, new_n12171,
    new_n12172, new_n12173, new_n12174, new_n12175, new_n12176, new_n12177,
    new_n12178, new_n12179, new_n12180, new_n12181, new_n12182, new_n12183,
    new_n12184, new_n12185, new_n12186, new_n12187, new_n12188, new_n12189,
    new_n12191, new_n12192, new_n12193, new_n12194, new_n12195, new_n12196,
    new_n12197, new_n12198, new_n12199, new_n12200, new_n12201, new_n12202,
    new_n12203, new_n12204, new_n12205, new_n12206, new_n12207, new_n12208,
    new_n12209, new_n12210, new_n12211, new_n12212, new_n12213, new_n12214,
    new_n12215, new_n12216, new_n12217, new_n12218, new_n12219, new_n12220,
    new_n12221, new_n12222, new_n12223, new_n12224, new_n12225, new_n12226,
    new_n12227, new_n12228, new_n12229, new_n12230, new_n12231, new_n12232,
    new_n12233, new_n12234, new_n12235, new_n12236, new_n12237, new_n12238,
    new_n12239, new_n12240, new_n12241, new_n12242, new_n12243, new_n12244,
    new_n12245, new_n12246, new_n12247, new_n12248, new_n12249, new_n12250,
    new_n12251, new_n12252, new_n12253, new_n12254, new_n12255, new_n12256,
    new_n12257, new_n12258, new_n12259, new_n12260, new_n12261, new_n12262,
    new_n12263, new_n12264, new_n12265, new_n12266, new_n12267, new_n12268,
    new_n12269, new_n12270, new_n12271, new_n12272, new_n12273, new_n12274,
    new_n12275, new_n12276, new_n12277, new_n12278, new_n12279, new_n12280,
    new_n12281, new_n12282, new_n12283, new_n12284, new_n12285, new_n12286,
    new_n12287, new_n12288, new_n12289, new_n12290, new_n12291, new_n12292,
    new_n12293, new_n12294, new_n12295, new_n12296, new_n12297, new_n12298,
    new_n12299, new_n12300, new_n12301, new_n12302, new_n12303, new_n12304,
    new_n12305, new_n12306, new_n12307, new_n12308, new_n12309, new_n12310,
    new_n12311, new_n12312, new_n12313, new_n12314, new_n12315, new_n12316,
    new_n12317, new_n12318, new_n12319, new_n12320, new_n12321, new_n12322,
    new_n12323, new_n12324, new_n12325, new_n12326, new_n12327, new_n12328,
    new_n12329, new_n12330, new_n12331, new_n12332, new_n12333, new_n12334,
    new_n12335, new_n12336, new_n12337, new_n12338, new_n12339, new_n12340,
    new_n12341, new_n12342, new_n12343, new_n12344, new_n12345, new_n12346,
    new_n12347, new_n12348, new_n12349, new_n12350, new_n12351, new_n12352,
    new_n12353, new_n12354, new_n12355, new_n12356, new_n12357, new_n12358,
    new_n12359, new_n12360, new_n12361, new_n12362, new_n12363, new_n12364,
    new_n12365, new_n12366, new_n12367, new_n12368, new_n12369, new_n12370,
    new_n12371, new_n12372, new_n12373, new_n12374, new_n12375, new_n12376,
    new_n12377, new_n12378, new_n12379, new_n12380, new_n12381, new_n12382,
    new_n12383, new_n12384, new_n12385, new_n12386, new_n12387, new_n12388,
    new_n12389, new_n12390, new_n12391, new_n12392, new_n12393, new_n12394,
    new_n12395, new_n12396, new_n12397, new_n12398, new_n12399, new_n12400,
    new_n12401, new_n12402, new_n12403, new_n12404, new_n12405, new_n12406,
    new_n12407, new_n12408, new_n12409, new_n12410, new_n12411, new_n12412,
    new_n12413, new_n12414, new_n12415, new_n12416, new_n12417, new_n12418,
    new_n12419, new_n12420, new_n12421, new_n12422, new_n12423, new_n12424,
    new_n12425, new_n12426, new_n12427, new_n12428, new_n12429, new_n12430,
    new_n12431, new_n12432, new_n12433, new_n12434, new_n12435, new_n12436,
    new_n12437, new_n12438, new_n12439, new_n12440, new_n12441, new_n12442,
    new_n12443, new_n12444, new_n12445, new_n12446, new_n12447, new_n12448,
    new_n12449, new_n12450, new_n12451, new_n12452, new_n12453, new_n12454,
    new_n12455, new_n12456, new_n12457, new_n12458, new_n12459, new_n12460,
    new_n12461, new_n12462, new_n12463, new_n12464, new_n12465, new_n12466,
    new_n12467, new_n12468, new_n12469, new_n12470, new_n12471, new_n12472,
    new_n12473, new_n12474, new_n12475, new_n12476, new_n12477, new_n12478,
    new_n12479, new_n12480, new_n12481, new_n12482, new_n12483, new_n12484,
    new_n12485, new_n12486, new_n12487, new_n12488, new_n12489, new_n12490,
    new_n12491, new_n12492, new_n12493, new_n12494, new_n12495, new_n12496,
    new_n12497, new_n12498, new_n12499, new_n12500, new_n12501, new_n12502,
    new_n12503, new_n12504, new_n12505, new_n12506, new_n12507, new_n12508,
    new_n12509, new_n12510, new_n12511, new_n12512, new_n12513, new_n12514,
    new_n12515, new_n12516, new_n12517, new_n12518, new_n12519, new_n12520,
    new_n12521, new_n12522, new_n12523, new_n12524, new_n12525, new_n12526,
    new_n12527, new_n12528, new_n12529, new_n12530, new_n12531, new_n12532,
    new_n12533, new_n12534, new_n12535, new_n12536, new_n12537, new_n12538,
    new_n12539, new_n12540, new_n12541, new_n12542, new_n12543, new_n12544,
    new_n12545, new_n12546, new_n12547, new_n12548, new_n12549, new_n12550,
    new_n12552, new_n12553, new_n12554, new_n12555, new_n12556, new_n12557,
    new_n12558, new_n12559, new_n12560, new_n12561, new_n12562, new_n12563,
    new_n12564, new_n12565, new_n12566, new_n12567, new_n12568, new_n12569,
    new_n12570, new_n12571, new_n12572, new_n12573, new_n12574, new_n12575,
    new_n12576, new_n12577, new_n12578, new_n12579, new_n12580, new_n12581,
    new_n12582, new_n12583, new_n12584, new_n12585, new_n12586, new_n12587,
    new_n12588, new_n12589, new_n12590, new_n12591, new_n12592, new_n12593,
    new_n12594, new_n12595, new_n12596, new_n12597, new_n12598, new_n12599,
    new_n12600, new_n12601, new_n12602, new_n12603, new_n12604, new_n12605,
    new_n12606, new_n12607, new_n12608, new_n12609, new_n12610, new_n12611,
    new_n12612, new_n12613, new_n12614, new_n12615, new_n12616, new_n12617,
    new_n12618, new_n12619, new_n12620, new_n12621, new_n12622, new_n12623,
    new_n12624, new_n12625, new_n12626, new_n12627, new_n12628, new_n12629,
    new_n12630, new_n12631, new_n12632, new_n12633, new_n12634, new_n12635,
    new_n12636, new_n12637, new_n12638, new_n12639, new_n12640, new_n12641,
    new_n12642, new_n12643, new_n12644, new_n12645, new_n12646, new_n12647,
    new_n12648, new_n12649, new_n12650, new_n12651, new_n12652, new_n12653,
    new_n12654, new_n12655, new_n12656, new_n12657, new_n12658, new_n12659,
    new_n12660, new_n12661, new_n12662, new_n12663, new_n12664, new_n12665,
    new_n12666, new_n12667, new_n12668, new_n12669, new_n12670, new_n12671,
    new_n12672, new_n12673, new_n12674, new_n12675, new_n12676, new_n12677,
    new_n12678, new_n12679, new_n12680, new_n12681, new_n12682, new_n12683,
    new_n12684, new_n12685, new_n12686, new_n12687, new_n12688, new_n12689,
    new_n12690, new_n12691, new_n12692, new_n12693, new_n12694, new_n12695,
    new_n12696, new_n12697, new_n12698, new_n12699, new_n12700, new_n12701,
    new_n12702, new_n12703, new_n12704, new_n12705, new_n12706, new_n12707,
    new_n12708, new_n12709, new_n12710, new_n12711, new_n12712, new_n12713,
    new_n12714, new_n12715, new_n12716, new_n12717, new_n12718, new_n12719,
    new_n12720, new_n12721, new_n12722, new_n12723, new_n12724, new_n12725,
    new_n12726, new_n12727, new_n12728, new_n12729, new_n12730, new_n12731,
    new_n12732, new_n12733, new_n12734, new_n12735, new_n12736, new_n12737,
    new_n12738, new_n12739, new_n12740, new_n12741, new_n12742, new_n12743,
    new_n12744, new_n12745, new_n12746, new_n12747, new_n12748, new_n12749,
    new_n12750, new_n12751, new_n12752, new_n12753, new_n12754, new_n12755,
    new_n12756, new_n12757, new_n12758, new_n12759, new_n12760, new_n12761,
    new_n12762, new_n12763, new_n12764, new_n12765, new_n12766, new_n12767,
    new_n12768, new_n12769, new_n12770, new_n12771, new_n12772, new_n12773,
    new_n12774, new_n12775, new_n12776, new_n12777, new_n12778, new_n12779,
    new_n12780, new_n12781, new_n12782, new_n12783, new_n12784, new_n12785,
    new_n12786, new_n12787, new_n12788, new_n12789, new_n12790, new_n12791,
    new_n12792, new_n12793, new_n12794, new_n12795, new_n12796, new_n12797,
    new_n12798, new_n12799, new_n12800, new_n12801, new_n12802, new_n12803,
    new_n12804, new_n12805, new_n12806, new_n12807, new_n12808, new_n12809,
    new_n12810, new_n12811, new_n12812, new_n12813, new_n12814, new_n12815,
    new_n12816, new_n12817, new_n12818, new_n12819, new_n12820, new_n12821,
    new_n12822, new_n12823, new_n12824, new_n12825, new_n12826, new_n12827,
    new_n12828, new_n12829, new_n12830, new_n12831, new_n12832, new_n12833,
    new_n12834, new_n12835, new_n12836, new_n12837, new_n12838, new_n12839,
    new_n12840, new_n12841, new_n12842, new_n12843, new_n12844, new_n12845,
    new_n12846, new_n12847, new_n12848, new_n12849, new_n12850, new_n12851,
    new_n12852, new_n12853, new_n12854, new_n12855, new_n12856, new_n12857,
    new_n12858, new_n12859, new_n12860, new_n12861, new_n12862, new_n12863,
    new_n12864, new_n12865, new_n12866, new_n12867, new_n12868, new_n12869,
    new_n12870, new_n12871, new_n12872, new_n12873, new_n12874, new_n12875,
    new_n12876, new_n12877, new_n12878, new_n12879, new_n12880, new_n12881,
    new_n12882, new_n12883, new_n12884, new_n12885, new_n12886, new_n12887,
    new_n12888, new_n12889, new_n12890, new_n12891, new_n12892, new_n12893,
    new_n12894, new_n12895, new_n12896, new_n12897, new_n12898, new_n12899,
    new_n12900, new_n12901, new_n12902, new_n12903, new_n12904, new_n12905,
    new_n12906, new_n12907, new_n12909, new_n12910, new_n12911, new_n12912,
    new_n12913, new_n12914, new_n12915, new_n12916, new_n12917, new_n12918,
    new_n12919, new_n12920, new_n12921, new_n12922, new_n12923, new_n12924,
    new_n12925, new_n12926, new_n12927, new_n12928, new_n12929, new_n12930,
    new_n12931, new_n12932, new_n12933, new_n12934, new_n12935, new_n12936,
    new_n12937, new_n12938, new_n12939, new_n12940, new_n12941, new_n12942,
    new_n12943, new_n12944, new_n12945, new_n12946, new_n12947, new_n12948,
    new_n12949, new_n12950, new_n12951, new_n12952, new_n12953, new_n12954,
    new_n12955, new_n12956, new_n12957, new_n12958, new_n12959, new_n12960,
    new_n12961, new_n12962, new_n12963, new_n12964, new_n12965, new_n12966,
    new_n12967, new_n12968, new_n12969, new_n12970, new_n12971, new_n12972,
    new_n12973, new_n12974, new_n12975, new_n12976, new_n12977, new_n12978,
    new_n12979, new_n12980, new_n12981, new_n12982, new_n12983, new_n12984,
    new_n12985, new_n12986, new_n12987, new_n12988, new_n12989, new_n12990,
    new_n12991, new_n12992, new_n12993, new_n12994, new_n12995, new_n12996,
    new_n12997, new_n12998, new_n12999, new_n13000, new_n13001, new_n13002,
    new_n13003, new_n13004, new_n13005, new_n13006, new_n13007, new_n13008,
    new_n13009, new_n13010, new_n13011, new_n13012, new_n13013, new_n13014,
    new_n13015, new_n13016, new_n13017, new_n13018, new_n13019, new_n13020,
    new_n13021, new_n13022, new_n13023, new_n13024, new_n13025, new_n13026,
    new_n13027, new_n13028, new_n13029, new_n13030, new_n13031, new_n13032,
    new_n13033, new_n13034, new_n13035, new_n13036, new_n13037, new_n13038,
    new_n13039, new_n13040, new_n13041, new_n13042, new_n13043, new_n13044,
    new_n13045, new_n13046, new_n13047, new_n13048, new_n13049, new_n13050,
    new_n13051, new_n13052, new_n13053, new_n13054, new_n13055, new_n13056,
    new_n13057, new_n13058, new_n13059, new_n13060, new_n13061, new_n13062,
    new_n13063, new_n13064, new_n13065, new_n13066, new_n13067, new_n13068,
    new_n13069, new_n13070, new_n13071, new_n13072, new_n13073, new_n13074,
    new_n13075, new_n13076, new_n13077, new_n13078, new_n13079, new_n13080,
    new_n13081, new_n13082, new_n13083, new_n13084, new_n13085, new_n13086,
    new_n13087, new_n13088, new_n13089, new_n13090, new_n13091, new_n13092,
    new_n13093, new_n13094, new_n13095, new_n13096, new_n13097, new_n13098,
    new_n13099, new_n13100, new_n13101, new_n13102, new_n13103, new_n13104,
    new_n13105, new_n13106, new_n13107, new_n13108, new_n13109, new_n13110,
    new_n13111, new_n13112, new_n13113, new_n13114, new_n13115, new_n13116,
    new_n13117, new_n13118, new_n13119, new_n13120, new_n13121, new_n13122,
    new_n13123, new_n13124, new_n13125, new_n13126, new_n13127, new_n13128,
    new_n13129, new_n13130, new_n13131, new_n13132, new_n13133, new_n13134,
    new_n13135, new_n13136, new_n13137, new_n13138, new_n13139, new_n13140,
    new_n13141, new_n13142, new_n13143, new_n13144, new_n13145, new_n13146,
    new_n13147, new_n13148, new_n13149, new_n13150, new_n13151, new_n13152,
    new_n13153, new_n13154, new_n13155, new_n13156, new_n13157, new_n13158,
    new_n13159, new_n13160, new_n13161, new_n13162, new_n13163, new_n13164,
    new_n13165, new_n13166, new_n13167, new_n13168, new_n13169, new_n13170,
    new_n13171, new_n13172, new_n13173, new_n13174, new_n13175, new_n13176,
    new_n13177, new_n13178, new_n13179, new_n13180, new_n13181, new_n13182,
    new_n13183, new_n13184, new_n13185, new_n13186, new_n13187, new_n13188,
    new_n13189, new_n13190, new_n13191, new_n13192, new_n13193, new_n13194,
    new_n13195, new_n13196, new_n13197, new_n13198, new_n13199, new_n13200,
    new_n13201, new_n13202, new_n13203, new_n13204, new_n13205, new_n13206,
    new_n13207, new_n13208, new_n13209, new_n13210, new_n13211, new_n13212,
    new_n13213, new_n13214, new_n13215, new_n13216, new_n13217, new_n13218,
    new_n13219, new_n13220, new_n13221, new_n13222, new_n13223, new_n13224,
    new_n13225, new_n13226, new_n13227, new_n13228, new_n13229, new_n13230,
    new_n13231, new_n13232, new_n13233, new_n13234, new_n13235, new_n13236,
    new_n13237, new_n13238, new_n13239, new_n13240, new_n13241, new_n13242,
    new_n13243, new_n13244, new_n13245, new_n13246, new_n13247, new_n13248,
    new_n13249, new_n13250, new_n13251, new_n13252, new_n13253, new_n13254,
    new_n13256, new_n13257, new_n13258, new_n13259, new_n13260, new_n13261,
    new_n13262, new_n13263, new_n13264, new_n13265, new_n13266, new_n13267,
    new_n13268, new_n13269, new_n13270, new_n13271, new_n13272, new_n13273,
    new_n13274, new_n13275, new_n13276, new_n13277, new_n13278, new_n13279,
    new_n13280, new_n13281, new_n13282, new_n13283, new_n13284, new_n13285,
    new_n13286, new_n13287, new_n13288, new_n13289, new_n13290, new_n13291,
    new_n13292, new_n13293, new_n13294, new_n13295, new_n13296, new_n13297,
    new_n13298, new_n13299, new_n13300, new_n13301, new_n13302, new_n13303,
    new_n13304, new_n13305, new_n13306, new_n13307, new_n13308, new_n13309,
    new_n13310, new_n13311, new_n13312, new_n13313, new_n13314, new_n13315,
    new_n13316, new_n13317, new_n13318, new_n13319, new_n13320, new_n13321,
    new_n13322, new_n13323, new_n13324, new_n13325, new_n13326, new_n13327,
    new_n13328, new_n13329, new_n13330, new_n13331, new_n13332, new_n13333,
    new_n13334, new_n13335, new_n13336, new_n13337, new_n13338, new_n13339,
    new_n13340, new_n13341, new_n13342, new_n13343, new_n13344, new_n13345,
    new_n13346, new_n13347, new_n13348, new_n13349, new_n13350, new_n13351,
    new_n13352, new_n13353, new_n13354, new_n13355, new_n13356, new_n13357,
    new_n13358, new_n13359, new_n13360, new_n13361, new_n13362, new_n13363,
    new_n13364, new_n13365, new_n13366, new_n13367, new_n13368, new_n13369,
    new_n13370, new_n13371, new_n13372, new_n13373, new_n13374, new_n13375,
    new_n13376, new_n13377, new_n13378, new_n13379, new_n13380, new_n13381,
    new_n13382, new_n13383, new_n13384, new_n13385, new_n13386, new_n13387,
    new_n13388, new_n13389, new_n13390, new_n13391, new_n13392, new_n13393,
    new_n13394, new_n13395, new_n13396, new_n13397, new_n13398, new_n13399,
    new_n13400, new_n13401, new_n13402, new_n13403, new_n13404, new_n13405,
    new_n13406, new_n13407, new_n13408, new_n13409, new_n13410, new_n13411,
    new_n13412, new_n13413, new_n13414, new_n13415, new_n13416, new_n13417,
    new_n13418, new_n13419, new_n13420, new_n13421, new_n13422, new_n13423,
    new_n13424, new_n13425, new_n13426, new_n13427, new_n13428, new_n13429,
    new_n13430, new_n13431, new_n13432, new_n13433, new_n13434, new_n13435,
    new_n13436, new_n13437, new_n13438, new_n13439, new_n13440, new_n13441,
    new_n13442, new_n13443, new_n13444, new_n13445, new_n13446, new_n13447,
    new_n13448, new_n13449, new_n13450, new_n13451, new_n13452, new_n13453,
    new_n13454, new_n13455, new_n13456, new_n13457, new_n13458, new_n13459,
    new_n13460, new_n13461, new_n13462, new_n13463, new_n13464, new_n13465,
    new_n13466, new_n13467, new_n13468, new_n13469, new_n13470, new_n13471,
    new_n13472, new_n13473, new_n13474, new_n13475, new_n13476, new_n13477,
    new_n13478, new_n13479, new_n13480, new_n13481, new_n13482, new_n13483,
    new_n13484, new_n13485, new_n13486, new_n13487, new_n13488, new_n13489,
    new_n13490, new_n13491, new_n13492, new_n13493, new_n13494, new_n13495,
    new_n13496, new_n13497, new_n13498, new_n13499, new_n13500, new_n13501,
    new_n13502, new_n13503, new_n13504, new_n13505, new_n13506, new_n13507,
    new_n13508, new_n13509, new_n13510, new_n13511, new_n13512, new_n13513,
    new_n13514, new_n13515, new_n13516, new_n13517, new_n13518, new_n13519,
    new_n13520, new_n13521, new_n13522, new_n13523, new_n13524, new_n13525,
    new_n13526, new_n13527, new_n13528, new_n13529, new_n13530, new_n13531,
    new_n13532, new_n13533, new_n13534, new_n13535, new_n13536, new_n13537,
    new_n13538, new_n13539, new_n13540, new_n13541, new_n13542, new_n13543,
    new_n13544, new_n13545, new_n13546, new_n13547, new_n13548, new_n13549,
    new_n13550, new_n13551, new_n13552, new_n13553, new_n13554, new_n13555,
    new_n13556, new_n13557, new_n13558, new_n13559, new_n13560, new_n13561,
    new_n13562, new_n13563, new_n13564, new_n13565, new_n13566, new_n13567,
    new_n13568, new_n13569, new_n13570, new_n13571, new_n13572, new_n13573,
    new_n13574, new_n13575, new_n13576, new_n13577, new_n13578, new_n13579,
    new_n13580, new_n13581, new_n13582, new_n13583, new_n13584, new_n13585,
    new_n13586, new_n13587, new_n13588, new_n13589, new_n13590, new_n13592,
    new_n13593, new_n13594, new_n13595, new_n13596, new_n13597, new_n13598,
    new_n13599, new_n13600, new_n13601, new_n13602, new_n13603, new_n13604,
    new_n13605, new_n13606, new_n13607, new_n13608, new_n13609, new_n13610,
    new_n13611, new_n13612, new_n13613, new_n13614, new_n13615, new_n13616,
    new_n13617, new_n13618, new_n13619, new_n13620, new_n13621, new_n13622,
    new_n13623, new_n13624, new_n13625, new_n13626, new_n13627, new_n13628,
    new_n13629, new_n13630, new_n13631, new_n13632, new_n13633, new_n13634,
    new_n13635, new_n13636, new_n13637, new_n13638, new_n13639, new_n13640,
    new_n13641, new_n13642, new_n13643, new_n13644, new_n13645, new_n13646,
    new_n13647, new_n13648, new_n13649, new_n13650, new_n13651, new_n13652,
    new_n13653, new_n13654, new_n13655, new_n13656, new_n13657, new_n13658,
    new_n13659, new_n13660, new_n13661, new_n13662, new_n13663, new_n13664,
    new_n13665, new_n13666, new_n13667, new_n13668, new_n13669, new_n13670,
    new_n13671, new_n13672, new_n13673, new_n13674, new_n13675, new_n13676,
    new_n13677, new_n13678, new_n13679, new_n13680, new_n13681, new_n13682,
    new_n13683, new_n13684, new_n13685, new_n13686, new_n13687, new_n13688,
    new_n13689, new_n13690, new_n13691, new_n13692, new_n13693, new_n13694,
    new_n13695, new_n13696, new_n13697, new_n13698, new_n13699, new_n13700,
    new_n13701, new_n13702, new_n13703, new_n13704, new_n13705, new_n13706,
    new_n13707, new_n13708, new_n13709, new_n13710, new_n13711, new_n13712,
    new_n13713, new_n13714, new_n13715, new_n13716, new_n13717, new_n13718,
    new_n13719, new_n13720, new_n13721, new_n13722, new_n13723, new_n13724,
    new_n13725, new_n13726, new_n13727, new_n13728, new_n13729, new_n13730,
    new_n13731, new_n13732, new_n13733, new_n13734, new_n13735, new_n13736,
    new_n13737, new_n13738, new_n13739, new_n13740, new_n13741, new_n13742,
    new_n13743, new_n13744, new_n13745, new_n13746, new_n13747, new_n13748,
    new_n13749, new_n13750, new_n13751, new_n13752, new_n13753, new_n13754,
    new_n13755, new_n13756, new_n13757, new_n13758, new_n13759, new_n13760,
    new_n13761, new_n13762, new_n13763, new_n13764, new_n13765, new_n13766,
    new_n13767, new_n13768, new_n13769, new_n13770, new_n13771, new_n13772,
    new_n13773, new_n13774, new_n13775, new_n13776, new_n13777, new_n13778,
    new_n13779, new_n13780, new_n13781, new_n13782, new_n13783, new_n13784,
    new_n13785, new_n13786, new_n13787, new_n13788, new_n13789, new_n13790,
    new_n13791, new_n13792, new_n13793, new_n13794, new_n13795, new_n13796,
    new_n13797, new_n13798, new_n13799, new_n13800, new_n13801, new_n13802,
    new_n13803, new_n13804, new_n13805, new_n13806, new_n13807, new_n13808,
    new_n13809, new_n13810, new_n13811, new_n13812, new_n13813, new_n13814,
    new_n13815, new_n13816, new_n13817, new_n13818, new_n13819, new_n13820,
    new_n13821, new_n13822, new_n13823, new_n13824, new_n13825, new_n13826,
    new_n13827, new_n13828, new_n13829, new_n13830, new_n13831, new_n13832,
    new_n13833, new_n13834, new_n13835, new_n13836, new_n13837, new_n13838,
    new_n13839, new_n13840, new_n13841, new_n13842, new_n13843, new_n13844,
    new_n13845, new_n13846, new_n13847, new_n13848, new_n13849, new_n13850,
    new_n13851, new_n13852, new_n13853, new_n13854, new_n13855, new_n13856,
    new_n13857, new_n13858, new_n13859, new_n13860, new_n13861, new_n13862,
    new_n13863, new_n13864, new_n13865, new_n13866, new_n13867, new_n13868,
    new_n13869, new_n13870, new_n13871, new_n13872, new_n13873, new_n13874,
    new_n13875, new_n13876, new_n13877, new_n13878, new_n13879, new_n13880,
    new_n13881, new_n13882, new_n13883, new_n13884, new_n13885, new_n13886,
    new_n13887, new_n13888, new_n13889, new_n13890, new_n13891, new_n13892,
    new_n13893, new_n13894, new_n13895, new_n13896, new_n13897, new_n13898,
    new_n13899, new_n13900, new_n13901, new_n13902, new_n13903, new_n13904,
    new_n13905, new_n13906, new_n13907, new_n13908, new_n13909, new_n13910,
    new_n13911, new_n13912, new_n13913, new_n13914, new_n13915, new_n13916,
    new_n13917, new_n13918, new_n13920, new_n13921, new_n13922, new_n13923,
    new_n13924, new_n13925, new_n13926, new_n13927, new_n13928, new_n13929,
    new_n13930, new_n13931, new_n13932, new_n13933, new_n13934, new_n13935,
    new_n13936, new_n13937, new_n13938, new_n13939, new_n13940, new_n13941,
    new_n13942, new_n13943, new_n13944, new_n13945, new_n13946, new_n13947,
    new_n13948, new_n13949, new_n13950, new_n13951, new_n13952, new_n13953,
    new_n13954, new_n13955, new_n13956, new_n13957, new_n13958, new_n13959,
    new_n13960, new_n13961, new_n13962, new_n13963, new_n13964, new_n13965,
    new_n13966, new_n13967, new_n13968, new_n13969, new_n13970, new_n13971,
    new_n13972, new_n13973, new_n13974, new_n13975, new_n13976, new_n13977,
    new_n13978, new_n13979, new_n13980, new_n13981, new_n13982, new_n13983,
    new_n13984, new_n13985, new_n13986, new_n13987, new_n13988, new_n13989,
    new_n13990, new_n13991, new_n13992, new_n13993, new_n13994, new_n13995,
    new_n13996, new_n13997, new_n13998, new_n13999, new_n14000, new_n14001,
    new_n14002, new_n14003, new_n14004, new_n14005, new_n14006, new_n14007,
    new_n14008, new_n14009, new_n14010, new_n14011, new_n14012, new_n14013,
    new_n14014, new_n14015, new_n14016, new_n14017, new_n14018, new_n14019,
    new_n14020, new_n14021, new_n14022, new_n14023, new_n14024, new_n14025,
    new_n14026, new_n14027, new_n14028, new_n14029, new_n14030, new_n14031,
    new_n14032, new_n14033, new_n14034, new_n14035, new_n14036, new_n14037,
    new_n14038, new_n14039, new_n14040, new_n14041, new_n14042, new_n14043,
    new_n14044, new_n14045, new_n14046, new_n14047, new_n14048, new_n14049,
    new_n14050, new_n14051, new_n14052, new_n14053, new_n14054, new_n14055,
    new_n14056, new_n14057, new_n14058, new_n14059, new_n14060, new_n14061,
    new_n14062, new_n14063, new_n14064, new_n14065, new_n14066, new_n14067,
    new_n14068, new_n14069, new_n14070, new_n14071, new_n14072, new_n14073,
    new_n14074, new_n14075, new_n14076, new_n14077, new_n14078, new_n14079,
    new_n14080, new_n14081, new_n14082, new_n14083, new_n14084, new_n14085,
    new_n14086, new_n14087, new_n14088, new_n14089, new_n14090, new_n14091,
    new_n14092, new_n14093, new_n14094, new_n14095, new_n14096, new_n14097,
    new_n14098, new_n14099, new_n14100, new_n14101, new_n14102, new_n14103,
    new_n14104, new_n14105, new_n14106, new_n14107, new_n14108, new_n14109,
    new_n14110, new_n14111, new_n14112, new_n14113, new_n14114, new_n14115,
    new_n14116, new_n14117, new_n14118, new_n14119, new_n14120, new_n14121,
    new_n14122, new_n14123, new_n14124, new_n14125, new_n14126, new_n14127,
    new_n14128, new_n14129, new_n14130, new_n14131, new_n14132, new_n14133,
    new_n14134, new_n14135, new_n14136, new_n14137, new_n14138, new_n14139,
    new_n14140, new_n14141, new_n14142, new_n14143, new_n14144, new_n14145,
    new_n14146, new_n14147, new_n14148, new_n14149, new_n14150, new_n14151,
    new_n14152, new_n14153, new_n14154, new_n14155, new_n14156, new_n14157,
    new_n14158, new_n14159, new_n14160, new_n14161, new_n14162, new_n14163,
    new_n14164, new_n14165, new_n14166, new_n14167, new_n14168, new_n14169,
    new_n14170, new_n14171, new_n14172, new_n14173, new_n14174, new_n14175,
    new_n14176, new_n14177, new_n14178, new_n14179, new_n14180, new_n14181,
    new_n14182, new_n14183, new_n14184, new_n14185, new_n14186, new_n14187,
    new_n14188, new_n14189, new_n14190, new_n14191, new_n14192, new_n14193,
    new_n14194, new_n14195, new_n14196, new_n14197, new_n14198, new_n14199,
    new_n14200, new_n14201, new_n14202, new_n14203, new_n14204, new_n14205,
    new_n14206, new_n14207, new_n14208, new_n14209, new_n14210, new_n14211,
    new_n14212, new_n14213, new_n14214, new_n14215, new_n14216, new_n14217,
    new_n14218, new_n14219, new_n14220, new_n14221, new_n14222, new_n14223,
    new_n14224, new_n14225, new_n14226, new_n14227, new_n14228, new_n14229,
    new_n14230, new_n14231, new_n14232, new_n14233, new_n14234, new_n14235,
    new_n14236, new_n14237, new_n14238, new_n14239, new_n14240, new_n14241,
    new_n14242, new_n14243, new_n14245, new_n14246, new_n14247, new_n14248,
    new_n14249, new_n14250, new_n14251, new_n14252, new_n14253, new_n14254,
    new_n14255, new_n14256, new_n14257, new_n14258, new_n14259, new_n14260,
    new_n14261, new_n14262, new_n14263, new_n14264, new_n14265, new_n14266,
    new_n14267, new_n14268, new_n14269, new_n14270, new_n14271, new_n14272,
    new_n14273, new_n14274, new_n14275, new_n14276, new_n14277, new_n14278,
    new_n14279, new_n14280, new_n14281, new_n14282, new_n14283, new_n14284,
    new_n14285, new_n14286, new_n14287, new_n14288, new_n14289, new_n14290,
    new_n14291, new_n14292, new_n14293, new_n14294, new_n14295, new_n14296,
    new_n14297, new_n14298, new_n14299, new_n14300, new_n14301, new_n14302,
    new_n14303, new_n14304, new_n14305, new_n14306, new_n14307, new_n14308,
    new_n14309, new_n14310, new_n14311, new_n14312, new_n14313, new_n14314,
    new_n14315, new_n14316, new_n14317, new_n14318, new_n14319, new_n14320,
    new_n14321, new_n14322, new_n14323, new_n14324, new_n14325, new_n14326,
    new_n14327, new_n14328, new_n14329, new_n14330, new_n14331, new_n14332,
    new_n14333, new_n14334, new_n14335, new_n14336, new_n14337, new_n14338,
    new_n14339, new_n14340, new_n14341, new_n14342, new_n14343, new_n14344,
    new_n14345, new_n14346, new_n14347, new_n14348, new_n14349, new_n14350,
    new_n14351, new_n14352, new_n14353, new_n14354, new_n14355, new_n14356,
    new_n14357, new_n14358, new_n14359, new_n14360, new_n14361, new_n14362,
    new_n14363, new_n14364, new_n14365, new_n14366, new_n14367, new_n14368,
    new_n14369, new_n14370, new_n14371, new_n14372, new_n14373, new_n14374,
    new_n14375, new_n14376, new_n14377, new_n14378, new_n14379, new_n14380,
    new_n14381, new_n14382, new_n14383, new_n14384, new_n14385, new_n14386,
    new_n14387, new_n14388, new_n14389, new_n14390, new_n14391, new_n14392,
    new_n14393, new_n14394, new_n14395, new_n14396, new_n14397, new_n14398,
    new_n14399, new_n14400, new_n14401, new_n14402, new_n14403, new_n14404,
    new_n14405, new_n14406, new_n14407, new_n14408, new_n14409, new_n14410,
    new_n14411, new_n14412, new_n14413, new_n14414, new_n14415, new_n14416,
    new_n14417, new_n14418, new_n14419, new_n14420, new_n14421, new_n14422,
    new_n14423, new_n14424, new_n14425, new_n14426, new_n14427, new_n14428,
    new_n14429, new_n14430, new_n14431, new_n14432, new_n14433, new_n14434,
    new_n14435, new_n14436, new_n14437, new_n14438, new_n14439, new_n14440,
    new_n14441, new_n14442, new_n14443, new_n14444, new_n14445, new_n14446,
    new_n14447, new_n14448, new_n14449, new_n14450, new_n14451, new_n14452,
    new_n14453, new_n14454, new_n14455, new_n14456, new_n14457, new_n14458,
    new_n14459, new_n14460, new_n14461, new_n14462, new_n14463, new_n14464,
    new_n14465, new_n14466, new_n14467, new_n14468, new_n14469, new_n14470,
    new_n14471, new_n14472, new_n14473, new_n14474, new_n14475, new_n14476,
    new_n14477, new_n14478, new_n14479, new_n14480, new_n14481, new_n14482,
    new_n14483, new_n14484, new_n14485, new_n14486, new_n14487, new_n14488,
    new_n14489, new_n14490, new_n14491, new_n14492, new_n14493, new_n14494,
    new_n14495, new_n14496, new_n14497, new_n14498, new_n14499, new_n14500,
    new_n14501, new_n14502, new_n14503, new_n14504, new_n14505, new_n14506,
    new_n14507, new_n14508, new_n14509, new_n14510, new_n14511, new_n14512,
    new_n14513, new_n14514, new_n14515, new_n14516, new_n14517, new_n14518,
    new_n14519, new_n14520, new_n14521, new_n14522, new_n14523, new_n14524,
    new_n14525, new_n14526, new_n14527, new_n14528, new_n14529, new_n14530,
    new_n14531, new_n14532, new_n14533, new_n14534, new_n14535, new_n14536,
    new_n14537, new_n14538, new_n14539, new_n14540, new_n14541, new_n14542,
    new_n14543, new_n14544, new_n14545, new_n14546, new_n14547, new_n14548,
    new_n14549, new_n14550, new_n14551, new_n14552, new_n14553, new_n14554,
    new_n14555, new_n14556, new_n14557, new_n14558, new_n14559, new_n14560,
    new_n14561, new_n14562, new_n14563, new_n14564, new_n14565, new_n14566,
    new_n14567, new_n14568, new_n14569, new_n14570, new_n14571, new_n14572,
    new_n14574, new_n14575, new_n14576, new_n14577, new_n14578, new_n14579,
    new_n14580, new_n14581, new_n14582, new_n14583, new_n14584, new_n14585,
    new_n14586, new_n14587, new_n14588, new_n14589, new_n14590, new_n14591,
    new_n14592, new_n14593, new_n14594, new_n14595, new_n14596, new_n14597,
    new_n14598, new_n14599, new_n14600, new_n14601, new_n14602, new_n14603,
    new_n14604, new_n14605, new_n14606, new_n14607, new_n14608, new_n14609,
    new_n14610, new_n14611, new_n14612, new_n14613, new_n14614, new_n14615,
    new_n14616, new_n14617, new_n14618, new_n14619, new_n14620, new_n14621,
    new_n14622, new_n14623, new_n14624, new_n14625, new_n14626, new_n14627,
    new_n14628, new_n14629, new_n14630, new_n14631, new_n14632, new_n14633,
    new_n14634, new_n14635, new_n14636, new_n14637, new_n14638, new_n14639,
    new_n14640, new_n14641, new_n14642, new_n14643, new_n14644, new_n14645,
    new_n14646, new_n14647, new_n14648, new_n14649, new_n14650, new_n14651,
    new_n14652, new_n14653, new_n14654, new_n14655, new_n14656, new_n14657,
    new_n14658, new_n14659, new_n14660, new_n14661, new_n14662, new_n14663,
    new_n14664, new_n14665, new_n14666, new_n14667, new_n14668, new_n14669,
    new_n14670, new_n14671, new_n14672, new_n14673, new_n14674, new_n14675,
    new_n14676, new_n14677, new_n14678, new_n14679, new_n14680, new_n14681,
    new_n14682, new_n14683, new_n14684, new_n14685, new_n14686, new_n14687,
    new_n14688, new_n14689, new_n14690, new_n14691, new_n14692, new_n14693,
    new_n14694, new_n14695, new_n14696, new_n14697, new_n14698, new_n14699,
    new_n14700, new_n14701, new_n14702, new_n14703, new_n14704, new_n14705,
    new_n14706, new_n14707, new_n14708, new_n14709, new_n14710, new_n14711,
    new_n14712, new_n14713, new_n14714, new_n14715, new_n14716, new_n14717,
    new_n14718, new_n14719, new_n14720, new_n14721, new_n14722, new_n14723,
    new_n14724, new_n14725, new_n14726, new_n14727, new_n14728, new_n14729,
    new_n14730, new_n14731, new_n14732, new_n14733, new_n14734, new_n14735,
    new_n14736, new_n14737, new_n14738, new_n14739, new_n14740, new_n14741,
    new_n14742, new_n14743, new_n14744, new_n14745, new_n14746, new_n14747,
    new_n14748, new_n14749, new_n14750, new_n14751, new_n14752, new_n14753,
    new_n14754, new_n14755, new_n14756, new_n14757, new_n14758, new_n14759,
    new_n14760, new_n14761, new_n14762, new_n14763, new_n14764, new_n14765,
    new_n14766, new_n14767, new_n14768, new_n14769, new_n14770, new_n14771,
    new_n14772, new_n14773, new_n14774, new_n14775, new_n14776, new_n14777,
    new_n14778, new_n14779, new_n14780, new_n14781, new_n14782, new_n14783,
    new_n14784, new_n14785, new_n14786, new_n14787, new_n14788, new_n14789,
    new_n14790, new_n14791, new_n14792, new_n14793, new_n14794, new_n14795,
    new_n14796, new_n14797, new_n14798, new_n14799, new_n14800, new_n14801,
    new_n14802, new_n14803, new_n14804, new_n14805, new_n14806, new_n14807,
    new_n14808, new_n14809, new_n14810, new_n14811, new_n14812, new_n14813,
    new_n14814, new_n14815, new_n14816, new_n14817, new_n14818, new_n14819,
    new_n14820, new_n14821, new_n14822, new_n14823, new_n14824, new_n14825,
    new_n14826, new_n14827, new_n14828, new_n14829, new_n14830, new_n14831,
    new_n14832, new_n14833, new_n14834, new_n14835, new_n14836, new_n14837,
    new_n14838, new_n14839, new_n14840, new_n14841, new_n14842, new_n14843,
    new_n14844, new_n14845, new_n14846, new_n14847, new_n14848, new_n14849,
    new_n14850, new_n14851, new_n14852, new_n14853, new_n14854, new_n14855,
    new_n14856, new_n14857, new_n14858, new_n14859, new_n14860, new_n14861,
    new_n14862, new_n14863, new_n14864, new_n14865, new_n14866, new_n14867,
    new_n14868, new_n14869, new_n14870, new_n14871, new_n14872, new_n14873,
    new_n14874, new_n14875, new_n14876, new_n14877, new_n14878, new_n14879,
    new_n14880, new_n14881, new_n14882, new_n14883, new_n14884, new_n14885,
    new_n14887, new_n14888, new_n14889, new_n14890, new_n14891, new_n14892,
    new_n14893, new_n14894, new_n14895, new_n14896, new_n14897, new_n14898,
    new_n14899, new_n14900, new_n14901, new_n14902, new_n14903, new_n14904,
    new_n14905, new_n14906, new_n14907, new_n14908, new_n14909, new_n14910,
    new_n14911, new_n14912, new_n14913, new_n14914, new_n14915, new_n14916,
    new_n14917, new_n14918, new_n14919, new_n14920, new_n14921, new_n14922,
    new_n14923, new_n14924, new_n14925, new_n14926, new_n14927, new_n14928,
    new_n14929, new_n14930, new_n14931, new_n14932, new_n14933, new_n14934,
    new_n14935, new_n14936, new_n14937, new_n14938, new_n14939, new_n14940,
    new_n14941, new_n14942, new_n14943, new_n14944, new_n14945, new_n14946,
    new_n14947, new_n14948, new_n14949, new_n14950, new_n14951, new_n14952,
    new_n14953, new_n14954, new_n14955, new_n14956, new_n14957, new_n14958,
    new_n14959, new_n14960, new_n14961, new_n14962, new_n14963, new_n14964,
    new_n14965, new_n14966, new_n14967, new_n14968, new_n14969, new_n14970,
    new_n14971, new_n14972, new_n14973, new_n14974, new_n14975, new_n14976,
    new_n14977, new_n14978, new_n14979, new_n14980, new_n14981, new_n14982,
    new_n14983, new_n14984, new_n14985, new_n14986, new_n14987, new_n14988,
    new_n14989, new_n14990, new_n14991, new_n14992, new_n14993, new_n14994,
    new_n14995, new_n14996, new_n14997, new_n14998, new_n14999, new_n15000,
    new_n15001, new_n15002, new_n15003, new_n15004, new_n15005, new_n15006,
    new_n15007, new_n15008, new_n15009, new_n15010, new_n15011, new_n15012,
    new_n15013, new_n15014, new_n15015, new_n15016, new_n15017, new_n15018,
    new_n15019, new_n15020, new_n15021, new_n15022, new_n15023, new_n15024,
    new_n15025, new_n15026, new_n15027, new_n15028, new_n15029, new_n15030,
    new_n15031, new_n15032, new_n15033, new_n15034, new_n15035, new_n15036,
    new_n15037, new_n15038, new_n15039, new_n15040, new_n15041, new_n15042,
    new_n15043, new_n15044, new_n15045, new_n15046, new_n15047, new_n15048,
    new_n15049, new_n15050, new_n15051, new_n15052, new_n15053, new_n15054,
    new_n15055, new_n15056, new_n15057, new_n15058, new_n15059, new_n15060,
    new_n15061, new_n15062, new_n15063, new_n15064, new_n15065, new_n15066,
    new_n15067, new_n15068, new_n15069, new_n15070, new_n15071, new_n15072,
    new_n15073, new_n15074, new_n15075, new_n15076, new_n15077, new_n15078,
    new_n15079, new_n15080, new_n15081, new_n15082, new_n15083, new_n15084,
    new_n15085, new_n15086, new_n15087, new_n15088, new_n15089, new_n15090,
    new_n15091, new_n15092, new_n15093, new_n15094, new_n15095, new_n15096,
    new_n15097, new_n15098, new_n15099, new_n15100, new_n15101, new_n15102,
    new_n15103, new_n15104, new_n15105, new_n15106, new_n15107, new_n15108,
    new_n15109, new_n15110, new_n15111, new_n15112, new_n15113, new_n15114,
    new_n15115, new_n15116, new_n15117, new_n15118, new_n15119, new_n15120,
    new_n15121, new_n15122, new_n15123, new_n15124, new_n15125, new_n15126,
    new_n15127, new_n15128, new_n15129, new_n15130, new_n15131, new_n15132,
    new_n15133, new_n15134, new_n15135, new_n15136, new_n15137, new_n15138,
    new_n15139, new_n15140, new_n15141, new_n15142, new_n15143, new_n15144,
    new_n15145, new_n15146, new_n15147, new_n15148, new_n15149, new_n15150,
    new_n15151, new_n15152, new_n15153, new_n15154, new_n15155, new_n15156,
    new_n15157, new_n15158, new_n15159, new_n15160, new_n15161, new_n15162,
    new_n15163, new_n15164, new_n15165, new_n15166, new_n15167, new_n15168,
    new_n15169, new_n15170, new_n15171, new_n15172, new_n15173, new_n15174,
    new_n15175, new_n15176, new_n15177, new_n15178, new_n15179, new_n15180,
    new_n15181, new_n15182, new_n15183, new_n15184, new_n15185, new_n15186,
    new_n15187, new_n15188, new_n15189, new_n15190, new_n15191, new_n15192,
    new_n15193, new_n15194, new_n15195, new_n15196, new_n15197, new_n15198,
    new_n15199, new_n15201, new_n15202, new_n15203, new_n15204, new_n15205,
    new_n15206, new_n15207, new_n15208, new_n15209, new_n15210, new_n15211,
    new_n15212, new_n15213, new_n15214, new_n15215, new_n15216, new_n15217,
    new_n15218, new_n15219, new_n15220, new_n15221, new_n15222, new_n15223,
    new_n15224, new_n15225, new_n15226, new_n15227, new_n15228, new_n15229,
    new_n15230, new_n15231, new_n15232, new_n15233, new_n15234, new_n15235,
    new_n15236, new_n15237, new_n15238, new_n15239, new_n15240, new_n15241,
    new_n15242, new_n15243, new_n15244, new_n15245, new_n15246, new_n15247,
    new_n15248, new_n15249, new_n15250, new_n15251, new_n15252, new_n15253,
    new_n15254, new_n15255, new_n15256, new_n15257, new_n15258, new_n15259,
    new_n15260, new_n15261, new_n15262, new_n15263, new_n15264, new_n15265,
    new_n15266, new_n15267, new_n15268, new_n15269, new_n15270, new_n15271,
    new_n15272, new_n15273, new_n15274, new_n15275, new_n15276, new_n15277,
    new_n15278, new_n15279, new_n15280, new_n15281, new_n15282, new_n15283,
    new_n15284, new_n15285, new_n15286, new_n15287, new_n15288, new_n15289,
    new_n15290, new_n15291, new_n15292, new_n15293, new_n15294, new_n15295,
    new_n15296, new_n15297, new_n15298, new_n15299, new_n15300, new_n15301,
    new_n15302, new_n15303, new_n15304, new_n15305, new_n15306, new_n15307,
    new_n15308, new_n15309, new_n15310, new_n15311, new_n15312, new_n15313,
    new_n15314, new_n15315, new_n15316, new_n15317, new_n15318, new_n15319,
    new_n15320, new_n15321, new_n15322, new_n15323, new_n15324, new_n15325,
    new_n15326, new_n15327, new_n15328, new_n15329, new_n15330, new_n15331,
    new_n15332, new_n15333, new_n15334, new_n15335, new_n15336, new_n15337,
    new_n15338, new_n15339, new_n15340, new_n15341, new_n15342, new_n15343,
    new_n15344, new_n15345, new_n15346, new_n15347, new_n15348, new_n15349,
    new_n15350, new_n15351, new_n15352, new_n15353, new_n15354, new_n15355,
    new_n15356, new_n15357, new_n15358, new_n15359, new_n15360, new_n15361,
    new_n15362, new_n15363, new_n15364, new_n15365, new_n15366, new_n15367,
    new_n15368, new_n15369, new_n15370, new_n15371, new_n15372, new_n15373,
    new_n15374, new_n15375, new_n15376, new_n15377, new_n15378, new_n15379,
    new_n15380, new_n15381, new_n15382, new_n15383, new_n15384, new_n15385,
    new_n15386, new_n15387, new_n15388, new_n15389, new_n15390, new_n15391,
    new_n15392, new_n15393, new_n15394, new_n15395, new_n15396, new_n15397,
    new_n15398, new_n15399, new_n15400, new_n15401, new_n15402, new_n15403,
    new_n15404, new_n15405, new_n15406, new_n15407, new_n15408, new_n15409,
    new_n15410, new_n15411, new_n15412, new_n15413, new_n15414, new_n15415,
    new_n15416, new_n15417, new_n15418, new_n15419, new_n15420, new_n15421,
    new_n15422, new_n15423, new_n15424, new_n15425, new_n15426, new_n15427,
    new_n15428, new_n15429, new_n15430, new_n15431, new_n15432, new_n15433,
    new_n15434, new_n15435, new_n15436, new_n15437, new_n15438, new_n15439,
    new_n15440, new_n15441, new_n15442, new_n15443, new_n15444, new_n15445,
    new_n15446, new_n15447, new_n15448, new_n15449, new_n15450, new_n15451,
    new_n15452, new_n15453, new_n15454, new_n15455, new_n15456, new_n15457,
    new_n15458, new_n15459, new_n15460, new_n15461, new_n15462, new_n15463,
    new_n15464, new_n15465, new_n15466, new_n15467, new_n15468, new_n15469,
    new_n15470, new_n15471, new_n15472, new_n15473, new_n15474, new_n15475,
    new_n15476, new_n15477, new_n15478, new_n15479, new_n15480, new_n15481,
    new_n15482, new_n15483, new_n15484, new_n15485, new_n15486, new_n15487,
    new_n15488, new_n15489, new_n15490, new_n15491, new_n15492, new_n15493,
    new_n15494, new_n15495, new_n15496, new_n15497, new_n15498, new_n15499,
    new_n15501, new_n15502, new_n15503, new_n15504, new_n15505, new_n15506,
    new_n15507, new_n15508, new_n15509, new_n15510, new_n15511, new_n15512,
    new_n15513, new_n15514, new_n15515, new_n15516, new_n15517, new_n15518,
    new_n15519, new_n15520, new_n15521, new_n15522, new_n15523, new_n15524,
    new_n15525, new_n15526, new_n15527, new_n15528, new_n15529, new_n15530,
    new_n15531, new_n15532, new_n15533, new_n15534, new_n15535, new_n15536,
    new_n15537, new_n15538, new_n15539, new_n15540, new_n15541, new_n15542,
    new_n15543, new_n15544, new_n15545, new_n15546, new_n15547, new_n15548,
    new_n15549, new_n15550, new_n15551, new_n15552, new_n15553, new_n15554,
    new_n15555, new_n15556, new_n15557, new_n15558, new_n15559, new_n15560,
    new_n15561, new_n15562, new_n15563, new_n15564, new_n15565, new_n15566,
    new_n15567, new_n15568, new_n15569, new_n15570, new_n15571, new_n15572,
    new_n15573, new_n15574, new_n15575, new_n15576, new_n15577, new_n15578,
    new_n15579, new_n15580, new_n15581, new_n15582, new_n15583, new_n15584,
    new_n15585, new_n15586, new_n15587, new_n15588, new_n15589, new_n15590,
    new_n15591, new_n15592, new_n15593, new_n15594, new_n15595, new_n15596,
    new_n15597, new_n15598, new_n15599, new_n15600, new_n15601, new_n15602,
    new_n15603, new_n15604, new_n15605, new_n15606, new_n15607, new_n15608,
    new_n15609, new_n15610, new_n15611, new_n15612, new_n15613, new_n15614,
    new_n15615, new_n15616, new_n15617, new_n15618, new_n15619, new_n15620,
    new_n15621, new_n15622, new_n15623, new_n15624, new_n15625, new_n15626,
    new_n15627, new_n15628, new_n15629, new_n15630, new_n15631, new_n15632,
    new_n15633, new_n15634, new_n15635, new_n15636, new_n15637, new_n15638,
    new_n15639, new_n15640, new_n15641, new_n15642, new_n15643, new_n15644,
    new_n15645, new_n15646, new_n15647, new_n15648, new_n15649, new_n15650,
    new_n15651, new_n15652, new_n15653, new_n15654, new_n15655, new_n15656,
    new_n15657, new_n15658, new_n15659, new_n15660, new_n15661, new_n15662,
    new_n15663, new_n15664, new_n15665, new_n15666, new_n15667, new_n15668,
    new_n15669, new_n15670, new_n15671, new_n15672, new_n15673, new_n15674,
    new_n15675, new_n15676, new_n15677, new_n15678, new_n15679, new_n15680,
    new_n15681, new_n15682, new_n15683, new_n15684, new_n15685, new_n15686,
    new_n15687, new_n15688, new_n15689, new_n15690, new_n15691, new_n15692,
    new_n15693, new_n15694, new_n15695, new_n15696, new_n15697, new_n15698,
    new_n15699, new_n15700, new_n15701, new_n15702, new_n15703, new_n15704,
    new_n15705, new_n15706, new_n15707, new_n15708, new_n15709, new_n15710,
    new_n15711, new_n15712, new_n15713, new_n15714, new_n15715, new_n15716,
    new_n15717, new_n15718, new_n15719, new_n15720, new_n15721, new_n15722,
    new_n15723, new_n15724, new_n15725, new_n15726, new_n15727, new_n15728,
    new_n15729, new_n15730, new_n15731, new_n15732, new_n15733, new_n15734,
    new_n15735, new_n15736, new_n15737, new_n15738, new_n15739, new_n15740,
    new_n15741, new_n15742, new_n15743, new_n15744, new_n15745, new_n15746,
    new_n15747, new_n15748, new_n15749, new_n15750, new_n15751, new_n15752,
    new_n15753, new_n15754, new_n15755, new_n15756, new_n15757, new_n15758,
    new_n15759, new_n15760, new_n15761, new_n15762, new_n15763, new_n15764,
    new_n15765, new_n15766, new_n15767, new_n15768, new_n15769, new_n15770,
    new_n15771, new_n15772, new_n15773, new_n15774, new_n15775, new_n15776,
    new_n15777, new_n15778, new_n15779, new_n15780, new_n15781, new_n15782,
    new_n15783, new_n15784, new_n15785, new_n15786, new_n15787, new_n15788,
    new_n15789, new_n15790, new_n15791, new_n15792, new_n15793, new_n15794,
    new_n15795, new_n15796, new_n15797, new_n15798, new_n15799, new_n15800,
    new_n15801, new_n15802, new_n15803, new_n15805, new_n15806, new_n15807,
    new_n15808, new_n15809, new_n15810, new_n15811, new_n15812, new_n15813,
    new_n15814, new_n15815, new_n15816, new_n15817, new_n15818, new_n15819,
    new_n15820, new_n15821, new_n15822, new_n15823, new_n15824, new_n15825,
    new_n15826, new_n15827, new_n15828, new_n15829, new_n15830, new_n15831,
    new_n15832, new_n15833, new_n15834, new_n15835, new_n15836, new_n15837,
    new_n15838, new_n15839, new_n15840, new_n15841, new_n15842, new_n15843,
    new_n15844, new_n15845, new_n15846, new_n15847, new_n15848, new_n15849,
    new_n15850, new_n15851, new_n15852, new_n15853, new_n15854, new_n15855,
    new_n15856, new_n15857, new_n15858, new_n15859, new_n15860, new_n15861,
    new_n15862, new_n15863, new_n15864, new_n15865, new_n15866, new_n15867,
    new_n15868, new_n15869, new_n15870, new_n15871, new_n15872, new_n15873,
    new_n15874, new_n15875, new_n15876, new_n15877, new_n15878, new_n15879,
    new_n15880, new_n15881, new_n15882, new_n15883, new_n15884, new_n15885,
    new_n15886, new_n15887, new_n15888, new_n15889, new_n15890, new_n15891,
    new_n15892, new_n15893, new_n15894, new_n15895, new_n15896, new_n15897,
    new_n15898, new_n15899, new_n15900, new_n15901, new_n15902, new_n15903,
    new_n15904, new_n15905, new_n15906, new_n15907, new_n15908, new_n15909,
    new_n15910, new_n15911, new_n15912, new_n15913, new_n15914, new_n15915,
    new_n15916, new_n15917, new_n15918, new_n15919, new_n15920, new_n15921,
    new_n15922, new_n15923, new_n15924, new_n15925, new_n15926, new_n15927,
    new_n15928, new_n15929, new_n15930, new_n15931, new_n15932, new_n15933,
    new_n15934, new_n15935, new_n15936, new_n15937, new_n15938, new_n15939,
    new_n15940, new_n15941, new_n15942, new_n15943, new_n15944, new_n15945,
    new_n15946, new_n15947, new_n15948, new_n15949, new_n15950, new_n15951,
    new_n15952, new_n15953, new_n15954, new_n15955, new_n15956, new_n15957,
    new_n15958, new_n15959, new_n15960, new_n15961, new_n15962, new_n15963,
    new_n15964, new_n15965, new_n15966, new_n15967, new_n15968, new_n15969,
    new_n15970, new_n15971, new_n15972, new_n15973, new_n15974, new_n15975,
    new_n15976, new_n15977, new_n15978, new_n15979, new_n15980, new_n15981,
    new_n15982, new_n15983, new_n15984, new_n15985, new_n15986, new_n15987,
    new_n15988, new_n15989, new_n15990, new_n15991, new_n15992, new_n15993,
    new_n15994, new_n15995, new_n15996, new_n15997, new_n15998, new_n15999,
    new_n16000, new_n16001, new_n16002, new_n16003, new_n16004, new_n16005,
    new_n16006, new_n16007, new_n16008, new_n16009, new_n16010, new_n16011,
    new_n16012, new_n16013, new_n16014, new_n16015, new_n16016, new_n16017,
    new_n16018, new_n16019, new_n16020, new_n16021, new_n16022, new_n16023,
    new_n16024, new_n16025, new_n16026, new_n16027, new_n16028, new_n16029,
    new_n16030, new_n16031, new_n16032, new_n16033, new_n16034, new_n16035,
    new_n16036, new_n16037, new_n16038, new_n16039, new_n16040, new_n16041,
    new_n16042, new_n16043, new_n16044, new_n16045, new_n16046, new_n16047,
    new_n16048, new_n16049, new_n16050, new_n16051, new_n16052, new_n16053,
    new_n16054, new_n16055, new_n16056, new_n16057, new_n16058, new_n16059,
    new_n16060, new_n16061, new_n16062, new_n16063, new_n16064, new_n16065,
    new_n16066, new_n16067, new_n16068, new_n16069, new_n16070, new_n16071,
    new_n16072, new_n16073, new_n16074, new_n16075, new_n16076, new_n16077,
    new_n16078, new_n16079, new_n16080, new_n16081, new_n16082, new_n16083,
    new_n16084, new_n16085, new_n16086, new_n16087, new_n16088, new_n16089,
    new_n16090, new_n16091, new_n16092, new_n16093, new_n16094, new_n16095,
    new_n16096, new_n16097, new_n16098, new_n16099, new_n16101, new_n16102,
    new_n16103, new_n16104, new_n16105, new_n16106, new_n16107, new_n16108,
    new_n16109, new_n16110, new_n16111, new_n16112, new_n16113, new_n16114,
    new_n16115, new_n16116, new_n16117, new_n16118, new_n16119, new_n16120,
    new_n16121, new_n16122, new_n16123, new_n16124, new_n16125, new_n16126,
    new_n16127, new_n16128, new_n16129, new_n16130, new_n16131, new_n16132,
    new_n16133, new_n16134, new_n16135, new_n16136, new_n16137, new_n16138,
    new_n16139, new_n16140, new_n16141, new_n16142, new_n16143, new_n16144,
    new_n16145, new_n16146, new_n16147, new_n16148, new_n16149, new_n16150,
    new_n16151, new_n16152, new_n16153, new_n16154, new_n16155, new_n16156,
    new_n16157, new_n16158, new_n16159, new_n16160, new_n16161, new_n16162,
    new_n16163, new_n16164, new_n16165, new_n16166, new_n16167, new_n16168,
    new_n16169, new_n16170, new_n16171, new_n16172, new_n16173, new_n16174,
    new_n16175, new_n16176, new_n16177, new_n16178, new_n16179, new_n16180,
    new_n16181, new_n16182, new_n16183, new_n16184, new_n16185, new_n16186,
    new_n16187, new_n16188, new_n16189, new_n16190, new_n16191, new_n16192,
    new_n16193, new_n16194, new_n16195, new_n16196, new_n16197, new_n16198,
    new_n16199, new_n16200, new_n16201, new_n16202, new_n16203, new_n16204,
    new_n16205, new_n16206, new_n16207, new_n16208, new_n16209, new_n16210,
    new_n16211, new_n16212, new_n16213, new_n16214, new_n16215, new_n16216,
    new_n16217, new_n16218, new_n16219, new_n16220, new_n16221, new_n16222,
    new_n16223, new_n16224, new_n16225, new_n16226, new_n16227, new_n16228,
    new_n16229, new_n16230, new_n16231, new_n16232, new_n16233, new_n16234,
    new_n16235, new_n16236, new_n16237, new_n16238, new_n16239, new_n16240,
    new_n16241, new_n16242, new_n16243, new_n16244, new_n16245, new_n16246,
    new_n16247, new_n16248, new_n16249, new_n16250, new_n16251, new_n16252,
    new_n16253, new_n16254, new_n16255, new_n16256, new_n16257, new_n16258,
    new_n16259, new_n16260, new_n16261, new_n16262, new_n16263, new_n16264,
    new_n16265, new_n16266, new_n16267, new_n16268, new_n16269, new_n16270,
    new_n16271, new_n16272, new_n16273, new_n16274, new_n16275, new_n16276,
    new_n16277, new_n16278, new_n16279, new_n16280, new_n16281, new_n16282,
    new_n16283, new_n16284, new_n16285, new_n16286, new_n16287, new_n16288,
    new_n16289, new_n16290, new_n16291, new_n16292, new_n16293, new_n16294,
    new_n16295, new_n16296, new_n16297, new_n16298, new_n16299, new_n16300,
    new_n16301, new_n16302, new_n16303, new_n16304, new_n16305, new_n16306,
    new_n16307, new_n16308, new_n16309, new_n16310, new_n16311, new_n16312,
    new_n16313, new_n16314, new_n16315, new_n16316, new_n16317, new_n16318,
    new_n16319, new_n16320, new_n16321, new_n16322, new_n16323, new_n16324,
    new_n16325, new_n16326, new_n16327, new_n16328, new_n16329, new_n16330,
    new_n16331, new_n16332, new_n16333, new_n16334, new_n16335, new_n16336,
    new_n16337, new_n16338, new_n16339, new_n16340, new_n16341, new_n16342,
    new_n16343, new_n16344, new_n16345, new_n16346, new_n16347, new_n16348,
    new_n16349, new_n16350, new_n16351, new_n16352, new_n16353, new_n16354,
    new_n16355, new_n16356, new_n16357, new_n16358, new_n16359, new_n16360,
    new_n16361, new_n16362, new_n16363, new_n16364, new_n16365, new_n16366,
    new_n16367, new_n16368, new_n16369, new_n16370, new_n16371, new_n16372,
    new_n16373, new_n16374, new_n16375, new_n16376, new_n16377, new_n16378,
    new_n16379, new_n16380, new_n16381, new_n16382, new_n16383, new_n16385,
    new_n16386, new_n16387, new_n16388, new_n16389, new_n16390, new_n16391,
    new_n16392, new_n16393, new_n16394, new_n16395, new_n16396, new_n16397,
    new_n16398, new_n16399, new_n16400, new_n16401, new_n16402, new_n16403,
    new_n16404, new_n16405, new_n16406, new_n16407, new_n16408, new_n16409,
    new_n16410, new_n16411, new_n16412, new_n16413, new_n16414, new_n16415,
    new_n16416, new_n16417, new_n16418, new_n16419, new_n16420, new_n16421,
    new_n16422, new_n16423, new_n16424, new_n16425, new_n16426, new_n16427,
    new_n16428, new_n16429, new_n16430, new_n16431, new_n16432, new_n16433,
    new_n16434, new_n16435, new_n16436, new_n16437, new_n16438, new_n16439,
    new_n16440, new_n16441, new_n16442, new_n16443, new_n16444, new_n16445,
    new_n16446, new_n16447, new_n16448, new_n16449, new_n16450, new_n16451,
    new_n16452, new_n16453, new_n16454, new_n16455, new_n16456, new_n16457,
    new_n16458, new_n16459, new_n16460, new_n16461, new_n16462, new_n16463,
    new_n16464, new_n16465, new_n16466, new_n16467, new_n16468, new_n16469,
    new_n16470, new_n16471, new_n16472, new_n16473, new_n16474, new_n16475,
    new_n16476, new_n16477, new_n16478, new_n16479, new_n16480, new_n16481,
    new_n16482, new_n16483, new_n16484, new_n16485, new_n16486, new_n16487,
    new_n16488, new_n16489, new_n16490, new_n16491, new_n16492, new_n16493,
    new_n16494, new_n16495, new_n16496, new_n16497, new_n16498, new_n16499,
    new_n16500, new_n16501, new_n16502, new_n16503, new_n16504, new_n16505,
    new_n16506, new_n16507, new_n16508, new_n16509, new_n16510, new_n16511,
    new_n16512, new_n16513, new_n16514, new_n16515, new_n16516, new_n16517,
    new_n16518, new_n16519, new_n16520, new_n16521, new_n16522, new_n16523,
    new_n16524, new_n16525, new_n16526, new_n16527, new_n16528, new_n16529,
    new_n16530, new_n16531, new_n16532, new_n16533, new_n16534, new_n16535,
    new_n16536, new_n16537, new_n16538, new_n16539, new_n16540, new_n16541,
    new_n16542, new_n16543, new_n16544, new_n16545, new_n16546, new_n16547,
    new_n16548, new_n16549, new_n16550, new_n16551, new_n16552, new_n16553,
    new_n16554, new_n16555, new_n16556, new_n16557, new_n16558, new_n16559,
    new_n16560, new_n16561, new_n16562, new_n16563, new_n16564, new_n16565,
    new_n16566, new_n16567, new_n16568, new_n16569, new_n16570, new_n16571,
    new_n16572, new_n16573, new_n16574, new_n16575, new_n16576, new_n16577,
    new_n16578, new_n16579, new_n16580, new_n16581, new_n16582, new_n16583,
    new_n16584, new_n16585, new_n16586, new_n16587, new_n16588, new_n16589,
    new_n16590, new_n16591, new_n16592, new_n16593, new_n16594, new_n16595,
    new_n16596, new_n16597, new_n16598, new_n16599, new_n16600, new_n16601,
    new_n16602, new_n16603, new_n16604, new_n16605, new_n16606, new_n16607,
    new_n16608, new_n16609, new_n16610, new_n16611, new_n16612, new_n16613,
    new_n16614, new_n16615, new_n16616, new_n16617, new_n16618, new_n16619,
    new_n16620, new_n16621, new_n16622, new_n16623, new_n16624, new_n16625,
    new_n16626, new_n16627, new_n16628, new_n16629, new_n16630, new_n16631,
    new_n16632, new_n16633, new_n16634, new_n16635, new_n16636, new_n16637,
    new_n16638, new_n16639, new_n16640, new_n16641, new_n16642, new_n16643,
    new_n16644, new_n16645, new_n16646, new_n16647, new_n16648, new_n16649,
    new_n16650, new_n16651, new_n16652, new_n16653, new_n16654, new_n16655,
    new_n16656, new_n16657, new_n16658, new_n16659, new_n16660, new_n16661,
    new_n16662, new_n16663, new_n16664, new_n16665, new_n16666, new_n16667,
    new_n16668, new_n16670, new_n16671, new_n16672, new_n16673, new_n16674,
    new_n16675, new_n16676, new_n16677, new_n16678, new_n16679, new_n16680,
    new_n16681, new_n16682, new_n16683, new_n16684, new_n16685, new_n16686,
    new_n16687, new_n16688, new_n16689, new_n16690, new_n16691, new_n16692,
    new_n16693, new_n16694, new_n16695, new_n16696, new_n16697, new_n16698,
    new_n16699, new_n16700, new_n16701, new_n16702, new_n16703, new_n16704,
    new_n16705, new_n16706, new_n16707, new_n16708, new_n16709, new_n16710,
    new_n16711, new_n16712, new_n16713, new_n16714, new_n16715, new_n16716,
    new_n16717, new_n16718, new_n16719, new_n16720, new_n16721, new_n16722,
    new_n16723, new_n16724, new_n16725, new_n16726, new_n16727, new_n16728,
    new_n16729, new_n16730, new_n16731, new_n16732, new_n16733, new_n16734,
    new_n16735, new_n16736, new_n16737, new_n16738, new_n16739, new_n16740,
    new_n16741, new_n16742, new_n16743, new_n16744, new_n16745, new_n16746,
    new_n16747, new_n16748, new_n16749, new_n16750, new_n16751, new_n16752,
    new_n16753, new_n16754, new_n16755, new_n16756, new_n16757, new_n16758,
    new_n16759, new_n16760, new_n16761, new_n16762, new_n16763, new_n16764,
    new_n16765, new_n16766, new_n16767, new_n16768, new_n16769, new_n16770,
    new_n16771, new_n16772, new_n16773, new_n16774, new_n16775, new_n16776,
    new_n16777, new_n16778, new_n16779, new_n16780, new_n16781, new_n16782,
    new_n16783, new_n16784, new_n16785, new_n16786, new_n16787, new_n16788,
    new_n16789, new_n16790, new_n16791, new_n16792, new_n16793, new_n16794,
    new_n16795, new_n16796, new_n16797, new_n16798, new_n16799, new_n16800,
    new_n16801, new_n16802, new_n16803, new_n16804, new_n16805, new_n16806,
    new_n16807, new_n16808, new_n16809, new_n16810, new_n16811, new_n16812,
    new_n16813, new_n16814, new_n16815, new_n16816, new_n16817, new_n16818,
    new_n16819, new_n16820, new_n16821, new_n16822, new_n16823, new_n16824,
    new_n16825, new_n16826, new_n16827, new_n16828, new_n16829, new_n16830,
    new_n16831, new_n16832, new_n16833, new_n16834, new_n16835, new_n16836,
    new_n16837, new_n16838, new_n16839, new_n16840, new_n16841, new_n16842,
    new_n16843, new_n16844, new_n16845, new_n16846, new_n16847, new_n16848,
    new_n16849, new_n16850, new_n16851, new_n16852, new_n16853, new_n16854,
    new_n16855, new_n16856, new_n16857, new_n16858, new_n16859, new_n16860,
    new_n16861, new_n16862, new_n16863, new_n16864, new_n16865, new_n16866,
    new_n16867, new_n16868, new_n16869, new_n16870, new_n16871, new_n16872,
    new_n16873, new_n16874, new_n16875, new_n16876, new_n16877, new_n16878,
    new_n16879, new_n16880, new_n16881, new_n16882, new_n16883, new_n16884,
    new_n16885, new_n16886, new_n16887, new_n16888, new_n16889, new_n16890,
    new_n16891, new_n16892, new_n16893, new_n16894, new_n16895, new_n16896,
    new_n16897, new_n16898, new_n16899, new_n16900, new_n16901, new_n16902,
    new_n16903, new_n16904, new_n16905, new_n16906, new_n16907, new_n16908,
    new_n16909, new_n16910, new_n16911, new_n16912, new_n16913, new_n16914,
    new_n16915, new_n16916, new_n16917, new_n16918, new_n16919, new_n16920,
    new_n16921, new_n16922, new_n16923, new_n16924, new_n16925, new_n16926,
    new_n16927, new_n16928, new_n16929, new_n16930, new_n16931, new_n16932,
    new_n16933, new_n16934, new_n16935, new_n16936, new_n16937, new_n16938,
    new_n16939, new_n16940, new_n16941, new_n16942, new_n16943, new_n16944,
    new_n16945, new_n16946, new_n16947, new_n16948, new_n16949, new_n16950,
    new_n16951, new_n16952, new_n16954, new_n16955, new_n16956, new_n16957,
    new_n16958, new_n16959, new_n16960, new_n16961, new_n16962, new_n16963,
    new_n16964, new_n16965, new_n16966, new_n16967, new_n16968, new_n16969,
    new_n16970, new_n16971, new_n16972, new_n16973, new_n16974, new_n16975,
    new_n16976, new_n16977, new_n16978, new_n16979, new_n16980, new_n16981,
    new_n16982, new_n16983, new_n16984, new_n16985, new_n16986, new_n16987,
    new_n16988, new_n16989, new_n16990, new_n16991, new_n16992, new_n16993,
    new_n16994, new_n16995, new_n16996, new_n16997, new_n16998, new_n16999,
    new_n17000, new_n17001, new_n17002, new_n17003, new_n17004, new_n17005,
    new_n17006, new_n17007, new_n17008, new_n17009, new_n17010, new_n17011,
    new_n17012, new_n17013, new_n17014, new_n17015, new_n17016, new_n17017,
    new_n17018, new_n17019, new_n17020, new_n17021, new_n17022, new_n17023,
    new_n17024, new_n17025, new_n17026, new_n17027, new_n17028, new_n17029,
    new_n17030, new_n17031, new_n17032, new_n17033, new_n17034, new_n17035,
    new_n17036, new_n17037, new_n17038, new_n17039, new_n17040, new_n17041,
    new_n17042, new_n17043, new_n17044, new_n17045, new_n17046, new_n17047,
    new_n17048, new_n17049, new_n17050, new_n17051, new_n17052, new_n17053,
    new_n17054, new_n17055, new_n17056, new_n17057, new_n17058, new_n17059,
    new_n17060, new_n17061, new_n17062, new_n17063, new_n17064, new_n17065,
    new_n17066, new_n17067, new_n17068, new_n17069, new_n17070, new_n17071,
    new_n17072, new_n17073, new_n17074, new_n17075, new_n17076, new_n17077,
    new_n17078, new_n17079, new_n17080, new_n17081, new_n17082, new_n17083,
    new_n17084, new_n17085, new_n17086, new_n17087, new_n17088, new_n17089,
    new_n17090, new_n17091, new_n17092, new_n17093, new_n17094, new_n17095,
    new_n17096, new_n17097, new_n17098, new_n17099, new_n17100, new_n17101,
    new_n17102, new_n17103, new_n17104, new_n17105, new_n17106, new_n17107,
    new_n17108, new_n17109, new_n17110, new_n17111, new_n17112, new_n17113,
    new_n17114, new_n17115, new_n17116, new_n17117, new_n17118, new_n17119,
    new_n17120, new_n17121, new_n17122, new_n17123, new_n17124, new_n17125,
    new_n17126, new_n17127, new_n17128, new_n17129, new_n17130, new_n17131,
    new_n17132, new_n17133, new_n17134, new_n17135, new_n17136, new_n17137,
    new_n17138, new_n17139, new_n17140, new_n17141, new_n17142, new_n17143,
    new_n17144, new_n17145, new_n17146, new_n17147, new_n17148, new_n17149,
    new_n17150, new_n17151, new_n17152, new_n17153, new_n17154, new_n17155,
    new_n17156, new_n17157, new_n17158, new_n17159, new_n17160, new_n17161,
    new_n17162, new_n17163, new_n17164, new_n17165, new_n17166, new_n17167,
    new_n17168, new_n17169, new_n17170, new_n17171, new_n17172, new_n17173,
    new_n17174, new_n17175, new_n17176, new_n17177, new_n17178, new_n17179,
    new_n17180, new_n17181, new_n17182, new_n17183, new_n17184, new_n17185,
    new_n17186, new_n17187, new_n17188, new_n17189, new_n17190, new_n17191,
    new_n17192, new_n17193, new_n17194, new_n17195, new_n17196, new_n17197,
    new_n17198, new_n17199, new_n17200, new_n17201, new_n17202, new_n17203,
    new_n17204, new_n17205, new_n17206, new_n17207, new_n17208, new_n17209,
    new_n17210, new_n17211, new_n17212, new_n17213, new_n17214, new_n17215,
    new_n17216, new_n17217, new_n17218, new_n17219, new_n17220, new_n17221,
    new_n17223, new_n17224, new_n17225, new_n17226, new_n17227, new_n17228,
    new_n17229, new_n17230, new_n17231, new_n17232, new_n17233, new_n17234,
    new_n17235, new_n17236, new_n17237, new_n17238, new_n17239, new_n17240,
    new_n17241, new_n17242, new_n17243, new_n17244, new_n17245, new_n17246,
    new_n17247, new_n17248, new_n17249, new_n17250, new_n17251, new_n17252,
    new_n17253, new_n17254, new_n17255, new_n17256, new_n17257, new_n17258,
    new_n17259, new_n17260, new_n17261, new_n17262, new_n17263, new_n17264,
    new_n17265, new_n17266, new_n17267, new_n17268, new_n17269, new_n17270,
    new_n17271, new_n17272, new_n17273, new_n17274, new_n17275, new_n17276,
    new_n17277, new_n17278, new_n17279, new_n17280, new_n17281, new_n17282,
    new_n17283, new_n17284, new_n17285, new_n17286, new_n17287, new_n17288,
    new_n17289, new_n17290, new_n17291, new_n17292, new_n17293, new_n17294,
    new_n17295, new_n17296, new_n17297, new_n17298, new_n17299, new_n17300,
    new_n17301, new_n17302, new_n17303, new_n17304, new_n17305, new_n17306,
    new_n17307, new_n17308, new_n17309, new_n17310, new_n17311, new_n17312,
    new_n17313, new_n17314, new_n17315, new_n17316, new_n17317, new_n17318,
    new_n17319, new_n17320, new_n17321, new_n17322, new_n17323, new_n17324,
    new_n17325, new_n17326, new_n17327, new_n17328, new_n17329, new_n17330,
    new_n17331, new_n17332, new_n17333, new_n17334, new_n17335, new_n17336,
    new_n17337, new_n17338, new_n17339, new_n17340, new_n17341, new_n17342,
    new_n17343, new_n17344, new_n17345, new_n17346, new_n17347, new_n17348,
    new_n17349, new_n17350, new_n17351, new_n17352, new_n17353, new_n17354,
    new_n17355, new_n17356, new_n17357, new_n17358, new_n17359, new_n17360,
    new_n17361, new_n17362, new_n17363, new_n17364, new_n17365, new_n17366,
    new_n17367, new_n17368, new_n17369, new_n17370, new_n17371, new_n17372,
    new_n17373, new_n17374, new_n17375, new_n17376, new_n17377, new_n17378,
    new_n17379, new_n17380, new_n17381, new_n17382, new_n17383, new_n17384,
    new_n17385, new_n17386, new_n17387, new_n17388, new_n17389, new_n17390,
    new_n17391, new_n17392, new_n17393, new_n17394, new_n17395, new_n17396,
    new_n17397, new_n17398, new_n17399, new_n17400, new_n17401, new_n17402,
    new_n17403, new_n17404, new_n17405, new_n17406, new_n17407, new_n17408,
    new_n17409, new_n17410, new_n17411, new_n17412, new_n17413, new_n17414,
    new_n17415, new_n17416, new_n17417, new_n17418, new_n17419, new_n17420,
    new_n17421, new_n17422, new_n17423, new_n17424, new_n17425, new_n17426,
    new_n17427, new_n17428, new_n17429, new_n17430, new_n17431, new_n17432,
    new_n17433, new_n17434, new_n17435, new_n17436, new_n17437, new_n17438,
    new_n17439, new_n17440, new_n17441, new_n17442, new_n17443, new_n17444,
    new_n17445, new_n17446, new_n17447, new_n17448, new_n17449, new_n17450,
    new_n17451, new_n17452, new_n17453, new_n17454, new_n17455, new_n17456,
    new_n17457, new_n17458, new_n17459, new_n17460, new_n17461, new_n17462,
    new_n17463, new_n17464, new_n17465, new_n17466, new_n17467, new_n17468,
    new_n17469, new_n17470, new_n17471, new_n17472, new_n17473, new_n17474,
    new_n17475, new_n17476, new_n17477, new_n17478, new_n17479, new_n17480,
    new_n17481, new_n17482, new_n17483, new_n17484, new_n17485, new_n17486,
    new_n17487, new_n17489, new_n17490, new_n17491, new_n17492, new_n17493,
    new_n17494, new_n17495, new_n17496, new_n17497, new_n17498, new_n17499,
    new_n17500, new_n17501, new_n17502, new_n17503, new_n17504, new_n17505,
    new_n17506, new_n17507, new_n17508, new_n17509, new_n17510, new_n17511,
    new_n17512, new_n17513, new_n17514, new_n17515, new_n17516, new_n17517,
    new_n17518, new_n17519, new_n17520, new_n17521, new_n17522, new_n17523,
    new_n17524, new_n17525, new_n17526, new_n17527, new_n17528, new_n17529,
    new_n17530, new_n17531, new_n17532, new_n17533, new_n17534, new_n17535,
    new_n17536, new_n17537, new_n17538, new_n17539, new_n17540, new_n17541,
    new_n17542, new_n17543, new_n17544, new_n17545, new_n17546, new_n17547,
    new_n17548, new_n17549, new_n17550, new_n17551, new_n17552, new_n17553,
    new_n17554, new_n17555, new_n17556, new_n17557, new_n17558, new_n17559,
    new_n17560, new_n17561, new_n17562, new_n17563, new_n17564, new_n17565,
    new_n17566, new_n17567, new_n17568, new_n17569, new_n17570, new_n17571,
    new_n17572, new_n17573, new_n17574, new_n17575, new_n17576, new_n17577,
    new_n17578, new_n17579, new_n17580, new_n17581, new_n17582, new_n17583,
    new_n17584, new_n17585, new_n17586, new_n17587, new_n17588, new_n17589,
    new_n17590, new_n17591, new_n17592, new_n17593, new_n17594, new_n17595,
    new_n17596, new_n17597, new_n17598, new_n17599, new_n17600, new_n17601,
    new_n17602, new_n17603, new_n17604, new_n17605, new_n17606, new_n17607,
    new_n17608, new_n17609, new_n17610, new_n17611, new_n17612, new_n17613,
    new_n17614, new_n17615, new_n17616, new_n17617, new_n17618, new_n17619,
    new_n17620, new_n17621, new_n17622, new_n17623, new_n17624, new_n17625,
    new_n17626, new_n17627, new_n17628, new_n17629, new_n17630, new_n17631,
    new_n17632, new_n17633, new_n17634, new_n17635, new_n17636, new_n17637,
    new_n17638, new_n17639, new_n17640, new_n17641, new_n17642, new_n17643,
    new_n17644, new_n17645, new_n17646, new_n17647, new_n17648, new_n17649,
    new_n17650, new_n17651, new_n17652, new_n17653, new_n17654, new_n17655,
    new_n17656, new_n17657, new_n17658, new_n17659, new_n17660, new_n17661,
    new_n17662, new_n17663, new_n17664, new_n17665, new_n17666, new_n17667,
    new_n17668, new_n17669, new_n17670, new_n17671, new_n17672, new_n17673,
    new_n17674, new_n17675, new_n17676, new_n17677, new_n17678, new_n17679,
    new_n17680, new_n17681, new_n17682, new_n17683, new_n17684, new_n17685,
    new_n17686, new_n17687, new_n17688, new_n17689, new_n17690, new_n17691,
    new_n17692, new_n17693, new_n17694, new_n17695, new_n17696, new_n17697,
    new_n17698, new_n17699, new_n17700, new_n17701, new_n17702, new_n17703,
    new_n17704, new_n17705, new_n17706, new_n17707, new_n17708, new_n17709,
    new_n17710, new_n17711, new_n17712, new_n17713, new_n17714, new_n17715,
    new_n17716, new_n17717, new_n17718, new_n17719, new_n17720, new_n17721,
    new_n17722, new_n17723, new_n17724, new_n17725, new_n17726, new_n17727,
    new_n17728, new_n17729, new_n17730, new_n17731, new_n17732, new_n17733,
    new_n17734, new_n17735, new_n17736, new_n17737, new_n17738, new_n17739,
    new_n17740, new_n17741, new_n17742, new_n17744, new_n17745, new_n17746,
    new_n17747, new_n17748, new_n17749, new_n17750, new_n17751, new_n17752,
    new_n17753, new_n17754, new_n17755, new_n17756, new_n17757, new_n17758,
    new_n17759, new_n17760, new_n17761, new_n17762, new_n17763, new_n17764,
    new_n17765, new_n17766, new_n17767, new_n17768, new_n17769, new_n17770,
    new_n17771, new_n17772, new_n17773, new_n17774, new_n17775, new_n17776,
    new_n17777, new_n17778, new_n17779, new_n17780, new_n17781, new_n17782,
    new_n17783, new_n17784, new_n17785, new_n17786, new_n17787, new_n17788,
    new_n17789, new_n17790, new_n17791, new_n17792, new_n17793, new_n17794,
    new_n17795, new_n17796, new_n17797, new_n17798, new_n17799, new_n17800,
    new_n17801, new_n17802, new_n17803, new_n17804, new_n17805, new_n17806,
    new_n17807, new_n17808, new_n17809, new_n17810, new_n17811, new_n17812,
    new_n17813, new_n17814, new_n17815, new_n17816, new_n17817, new_n17818,
    new_n17819, new_n17820, new_n17821, new_n17822, new_n17823, new_n17824,
    new_n17825, new_n17826, new_n17827, new_n17828, new_n17829, new_n17830,
    new_n17831, new_n17832, new_n17833, new_n17834, new_n17835, new_n17836,
    new_n17837, new_n17838, new_n17839, new_n17840, new_n17841, new_n17842,
    new_n17843, new_n17844, new_n17845, new_n17846, new_n17847, new_n17848,
    new_n17849, new_n17850, new_n17851, new_n17852, new_n17853, new_n17854,
    new_n17855, new_n17856, new_n17857, new_n17858, new_n17859, new_n17860,
    new_n17861, new_n17862, new_n17863, new_n17864, new_n17865, new_n17866,
    new_n17867, new_n17868, new_n17869, new_n17870, new_n17871, new_n17872,
    new_n17873, new_n17874, new_n17875, new_n17876, new_n17877, new_n17878,
    new_n17879, new_n17880, new_n17881, new_n17882, new_n17883, new_n17884,
    new_n17885, new_n17886, new_n17887, new_n17888, new_n17889, new_n17890,
    new_n17891, new_n17892, new_n17893, new_n17894, new_n17895, new_n17896,
    new_n17897, new_n17898, new_n17899, new_n17900, new_n17901, new_n17902,
    new_n17903, new_n17904, new_n17905, new_n17906, new_n17907, new_n17908,
    new_n17909, new_n17910, new_n17911, new_n17912, new_n17913, new_n17914,
    new_n17915, new_n17916, new_n17917, new_n17918, new_n17919, new_n17920,
    new_n17921, new_n17922, new_n17923, new_n17924, new_n17925, new_n17926,
    new_n17927, new_n17928, new_n17929, new_n17930, new_n17931, new_n17932,
    new_n17933, new_n17934, new_n17935, new_n17936, new_n17937, new_n17938,
    new_n17939, new_n17940, new_n17941, new_n17942, new_n17943, new_n17944,
    new_n17945, new_n17946, new_n17947, new_n17948, new_n17949, new_n17950,
    new_n17951, new_n17952, new_n17953, new_n17954, new_n17955, new_n17956,
    new_n17957, new_n17958, new_n17959, new_n17960, new_n17961, new_n17962,
    new_n17963, new_n17964, new_n17965, new_n17966, new_n17967, new_n17968,
    new_n17969, new_n17970, new_n17971, new_n17972, new_n17973, new_n17974,
    new_n17975, new_n17976, new_n17977, new_n17978, new_n17979, new_n17980,
    new_n17981, new_n17982, new_n17983, new_n17984, new_n17985, new_n17986,
    new_n17987, new_n17988, new_n17989, new_n17990, new_n17991, new_n17992,
    new_n17993, new_n17994, new_n17996, new_n17997, new_n17998, new_n17999,
    new_n18000, new_n18001, new_n18002, new_n18003, new_n18004, new_n18005,
    new_n18006, new_n18007, new_n18008, new_n18009, new_n18010, new_n18011,
    new_n18012, new_n18013, new_n18014, new_n18015, new_n18016, new_n18017,
    new_n18018, new_n18019, new_n18020, new_n18021, new_n18022, new_n18023,
    new_n18024, new_n18025, new_n18026, new_n18027, new_n18028, new_n18029,
    new_n18030, new_n18031, new_n18032, new_n18033, new_n18034, new_n18035,
    new_n18036, new_n18037, new_n18038, new_n18039, new_n18040, new_n18041,
    new_n18042, new_n18043, new_n18044, new_n18045, new_n18046, new_n18047,
    new_n18048, new_n18049, new_n18050, new_n18051, new_n18052, new_n18053,
    new_n18054, new_n18055, new_n18056, new_n18057, new_n18058, new_n18059,
    new_n18060, new_n18061, new_n18062, new_n18063, new_n18064, new_n18065,
    new_n18066, new_n18067, new_n18068, new_n18069, new_n18070, new_n18071,
    new_n18072, new_n18073, new_n18074, new_n18075, new_n18076, new_n18077,
    new_n18078, new_n18079, new_n18080, new_n18081, new_n18082, new_n18083,
    new_n18084, new_n18085, new_n18086, new_n18087, new_n18088, new_n18089,
    new_n18090, new_n18091, new_n18092, new_n18093, new_n18094, new_n18095,
    new_n18096, new_n18097, new_n18098, new_n18099, new_n18100, new_n18101,
    new_n18102, new_n18103, new_n18104, new_n18105, new_n18106, new_n18107,
    new_n18108, new_n18109, new_n18110, new_n18111, new_n18112, new_n18113,
    new_n18114, new_n18115, new_n18116, new_n18117, new_n18118, new_n18119,
    new_n18120, new_n18121, new_n18122, new_n18123, new_n18124, new_n18125,
    new_n18126, new_n18127, new_n18128, new_n18129, new_n18130, new_n18131,
    new_n18132, new_n18133, new_n18134, new_n18135, new_n18136, new_n18137,
    new_n18138, new_n18139, new_n18140, new_n18141, new_n18142, new_n18143,
    new_n18144, new_n18145, new_n18146, new_n18147, new_n18148, new_n18149,
    new_n18150, new_n18151, new_n18152, new_n18153, new_n18154, new_n18155,
    new_n18156, new_n18157, new_n18158, new_n18159, new_n18160, new_n18161,
    new_n18162, new_n18163, new_n18164, new_n18165, new_n18166, new_n18167,
    new_n18168, new_n18169, new_n18170, new_n18171, new_n18172, new_n18173,
    new_n18174, new_n18175, new_n18176, new_n18177, new_n18178, new_n18179,
    new_n18180, new_n18181, new_n18182, new_n18183, new_n18184, new_n18185,
    new_n18186, new_n18187, new_n18188, new_n18189, new_n18190, new_n18191,
    new_n18192, new_n18193, new_n18194, new_n18195, new_n18196, new_n18197,
    new_n18198, new_n18199, new_n18200, new_n18201, new_n18202, new_n18203,
    new_n18204, new_n18205, new_n18206, new_n18207, new_n18208, new_n18209,
    new_n18210, new_n18211, new_n18212, new_n18213, new_n18214, new_n18215,
    new_n18216, new_n18217, new_n18218, new_n18219, new_n18220, new_n18221,
    new_n18222, new_n18223, new_n18224, new_n18225, new_n18226, new_n18227,
    new_n18228, new_n18229, new_n18230, new_n18231, new_n18232, new_n18233,
    new_n18234, new_n18235, new_n18236, new_n18237, new_n18238, new_n18239,
    new_n18240, new_n18241, new_n18242, new_n18243, new_n18244, new_n18245,
    new_n18247, new_n18248, new_n18249, new_n18250, new_n18251, new_n18252,
    new_n18253, new_n18254, new_n18255, new_n18256, new_n18257, new_n18258,
    new_n18259, new_n18260, new_n18261, new_n18262, new_n18263, new_n18264,
    new_n18265, new_n18266, new_n18267, new_n18268, new_n18269, new_n18270,
    new_n18271, new_n18272, new_n18273, new_n18274, new_n18275, new_n18276,
    new_n18277, new_n18278, new_n18279, new_n18280, new_n18281, new_n18282,
    new_n18283, new_n18284, new_n18285, new_n18286, new_n18287, new_n18288,
    new_n18289, new_n18290, new_n18291, new_n18292, new_n18293, new_n18294,
    new_n18295, new_n18296, new_n18297, new_n18298, new_n18299, new_n18300,
    new_n18301, new_n18302, new_n18303, new_n18304, new_n18305, new_n18306,
    new_n18307, new_n18308, new_n18309, new_n18310, new_n18311, new_n18312,
    new_n18313, new_n18314, new_n18315, new_n18316, new_n18317, new_n18318,
    new_n18319, new_n18320, new_n18321, new_n18322, new_n18323, new_n18324,
    new_n18325, new_n18326, new_n18327, new_n18328, new_n18329, new_n18330,
    new_n18331, new_n18332, new_n18333, new_n18334, new_n18335, new_n18336,
    new_n18337, new_n18338, new_n18339, new_n18340, new_n18341, new_n18342,
    new_n18343, new_n18344, new_n18345, new_n18346, new_n18347, new_n18348,
    new_n18349, new_n18350, new_n18351, new_n18352, new_n18353, new_n18354,
    new_n18355, new_n18356, new_n18357, new_n18358, new_n18359, new_n18360,
    new_n18361, new_n18362, new_n18363, new_n18364, new_n18365, new_n18366,
    new_n18367, new_n18368, new_n18369, new_n18370, new_n18371, new_n18372,
    new_n18373, new_n18374, new_n18375, new_n18376, new_n18377, new_n18378,
    new_n18379, new_n18380, new_n18381, new_n18382, new_n18383, new_n18384,
    new_n18385, new_n18386, new_n18387, new_n18388, new_n18389, new_n18390,
    new_n18391, new_n18392, new_n18393, new_n18394, new_n18395, new_n18396,
    new_n18397, new_n18398, new_n18399, new_n18400, new_n18401, new_n18402,
    new_n18403, new_n18404, new_n18405, new_n18406, new_n18407, new_n18408,
    new_n18409, new_n18410, new_n18411, new_n18412, new_n18413, new_n18414,
    new_n18415, new_n18416, new_n18417, new_n18418, new_n18419, new_n18420,
    new_n18421, new_n18422, new_n18423, new_n18424, new_n18425, new_n18426,
    new_n18427, new_n18428, new_n18429, new_n18430, new_n18431, new_n18432,
    new_n18433, new_n18434, new_n18435, new_n18436, new_n18437, new_n18438,
    new_n18439, new_n18440, new_n18441, new_n18442, new_n18443, new_n18444,
    new_n18445, new_n18446, new_n18447, new_n18448, new_n18449, new_n18450,
    new_n18451, new_n18452, new_n18453, new_n18454, new_n18455, new_n18456,
    new_n18457, new_n18458, new_n18459, new_n18460, new_n18461, new_n18462,
    new_n18463, new_n18464, new_n18465, new_n18466, new_n18467, new_n18468,
    new_n18469, new_n18470, new_n18471, new_n18472, new_n18473, new_n18474,
    new_n18475, new_n18476, new_n18477, new_n18478, new_n18479, new_n18480,
    new_n18481, new_n18483, new_n18484, new_n18485, new_n18486, new_n18487,
    new_n18488, new_n18489, new_n18490, new_n18491, new_n18492, new_n18493,
    new_n18494, new_n18495, new_n18496, new_n18497, new_n18498, new_n18499,
    new_n18500, new_n18501, new_n18502, new_n18503, new_n18504, new_n18505,
    new_n18506, new_n18507, new_n18508, new_n18509, new_n18510, new_n18511,
    new_n18512, new_n18513, new_n18514, new_n18515, new_n18516, new_n18517,
    new_n18518, new_n18519, new_n18520, new_n18521, new_n18522, new_n18523,
    new_n18524, new_n18525, new_n18526, new_n18527, new_n18528, new_n18529,
    new_n18530, new_n18531, new_n18532, new_n18533, new_n18534, new_n18535,
    new_n18536, new_n18537, new_n18538, new_n18539, new_n18540, new_n18541,
    new_n18542, new_n18543, new_n18544, new_n18545, new_n18546, new_n18547,
    new_n18548, new_n18549, new_n18550, new_n18551, new_n18552, new_n18553,
    new_n18554, new_n18555, new_n18556, new_n18557, new_n18558, new_n18559,
    new_n18560, new_n18561, new_n18562, new_n18563, new_n18564, new_n18565,
    new_n18566, new_n18567, new_n18568, new_n18569, new_n18570, new_n18571,
    new_n18572, new_n18573, new_n18574, new_n18575, new_n18576, new_n18577,
    new_n18578, new_n18579, new_n18580, new_n18581, new_n18582, new_n18583,
    new_n18584, new_n18585, new_n18586, new_n18587, new_n18588, new_n18589,
    new_n18590, new_n18591, new_n18592, new_n18593, new_n18594, new_n18595,
    new_n18596, new_n18597, new_n18598, new_n18599, new_n18600, new_n18601,
    new_n18602, new_n18603, new_n18604, new_n18605, new_n18606, new_n18607,
    new_n18608, new_n18609, new_n18610, new_n18611, new_n18612, new_n18613,
    new_n18614, new_n18615, new_n18616, new_n18617, new_n18618, new_n18619,
    new_n18620, new_n18621, new_n18622, new_n18623, new_n18624, new_n18625,
    new_n18626, new_n18627, new_n18628, new_n18629, new_n18630, new_n18631,
    new_n18632, new_n18633, new_n18634, new_n18635, new_n18636, new_n18637,
    new_n18638, new_n18639, new_n18640, new_n18641, new_n18642, new_n18643,
    new_n18644, new_n18645, new_n18646, new_n18647, new_n18648, new_n18649,
    new_n18650, new_n18651, new_n18652, new_n18653, new_n18654, new_n18655,
    new_n18656, new_n18657, new_n18658, new_n18659, new_n18660, new_n18661,
    new_n18662, new_n18663, new_n18664, new_n18665, new_n18666, new_n18667,
    new_n18668, new_n18669, new_n18670, new_n18671, new_n18672, new_n18673,
    new_n18674, new_n18675, new_n18676, new_n18677, new_n18678, new_n18679,
    new_n18680, new_n18681, new_n18682, new_n18683, new_n18684, new_n18685,
    new_n18686, new_n18687, new_n18688, new_n18689, new_n18690, new_n18691,
    new_n18692, new_n18693, new_n18694, new_n18695, new_n18696, new_n18697,
    new_n18698, new_n18699, new_n18700, new_n18701, new_n18702, new_n18703,
    new_n18704, new_n18705, new_n18706, new_n18707, new_n18708, new_n18709,
    new_n18710, new_n18711, new_n18712, new_n18713, new_n18714, new_n18715,
    new_n18716, new_n18717, new_n18718, new_n18720, new_n18721, new_n18722,
    new_n18723, new_n18724, new_n18725, new_n18726, new_n18727, new_n18728,
    new_n18729, new_n18730, new_n18731, new_n18732, new_n18733, new_n18734,
    new_n18735, new_n18736, new_n18737, new_n18738, new_n18739, new_n18740,
    new_n18741, new_n18742, new_n18743, new_n18744, new_n18745, new_n18746,
    new_n18747, new_n18748, new_n18749, new_n18750, new_n18751, new_n18752,
    new_n18753, new_n18754, new_n18755, new_n18756, new_n18757, new_n18758,
    new_n18759, new_n18760, new_n18761, new_n18762, new_n18763, new_n18764,
    new_n18765, new_n18766, new_n18767, new_n18768, new_n18769, new_n18770,
    new_n18771, new_n18772, new_n18773, new_n18774, new_n18775, new_n18776,
    new_n18777, new_n18778, new_n18779, new_n18780, new_n18781, new_n18782,
    new_n18783, new_n18784, new_n18785, new_n18786, new_n18787, new_n18788,
    new_n18789, new_n18790, new_n18791, new_n18792, new_n18793, new_n18794,
    new_n18795, new_n18796, new_n18797, new_n18798, new_n18799, new_n18800,
    new_n18801, new_n18802, new_n18803, new_n18804, new_n18805, new_n18806,
    new_n18807, new_n18808, new_n18809, new_n18810, new_n18811, new_n18812,
    new_n18813, new_n18814, new_n18815, new_n18816, new_n18817, new_n18818,
    new_n18819, new_n18820, new_n18821, new_n18822, new_n18823, new_n18824,
    new_n18825, new_n18826, new_n18827, new_n18828, new_n18829, new_n18830,
    new_n18831, new_n18832, new_n18833, new_n18834, new_n18835, new_n18836,
    new_n18837, new_n18838, new_n18839, new_n18840, new_n18841, new_n18842,
    new_n18843, new_n18844, new_n18845, new_n18846, new_n18847, new_n18848,
    new_n18849, new_n18850, new_n18851, new_n18852, new_n18853, new_n18854,
    new_n18855, new_n18856, new_n18857, new_n18858, new_n18859, new_n18860,
    new_n18861, new_n18862, new_n18863, new_n18864, new_n18865, new_n18866,
    new_n18867, new_n18868, new_n18869, new_n18870, new_n18871, new_n18872,
    new_n18873, new_n18874, new_n18875, new_n18876, new_n18877, new_n18878,
    new_n18879, new_n18880, new_n18881, new_n18882, new_n18883, new_n18884,
    new_n18885, new_n18886, new_n18887, new_n18888, new_n18889, new_n18890,
    new_n18891, new_n18892, new_n18893, new_n18894, new_n18895, new_n18896,
    new_n18897, new_n18898, new_n18899, new_n18900, new_n18901, new_n18902,
    new_n18903, new_n18904, new_n18905, new_n18906, new_n18907, new_n18908,
    new_n18909, new_n18910, new_n18911, new_n18912, new_n18913, new_n18914,
    new_n18915, new_n18916, new_n18917, new_n18918, new_n18919, new_n18920,
    new_n18921, new_n18922, new_n18923, new_n18924, new_n18925, new_n18926,
    new_n18927, new_n18928, new_n18929, new_n18930, new_n18931, new_n18932,
    new_n18933, new_n18934, new_n18935, new_n18936, new_n18937, new_n18938,
    new_n18939, new_n18940, new_n18941, new_n18942, new_n18943, new_n18945,
    new_n18946, new_n18947, new_n18948, new_n18949, new_n18950, new_n18951,
    new_n18952, new_n18953, new_n18954, new_n18955, new_n18956, new_n18957,
    new_n18958, new_n18959, new_n18960, new_n18961, new_n18962, new_n18963,
    new_n18964, new_n18965, new_n18966, new_n18967, new_n18968, new_n18969,
    new_n18970, new_n18971, new_n18972, new_n18973, new_n18974, new_n18975,
    new_n18976, new_n18977, new_n18978, new_n18979, new_n18980, new_n18981,
    new_n18982, new_n18983, new_n18984, new_n18985, new_n18986, new_n18987,
    new_n18988, new_n18989, new_n18990, new_n18991, new_n18992, new_n18993,
    new_n18994, new_n18995, new_n18996, new_n18997, new_n18998, new_n18999,
    new_n19000, new_n19001, new_n19002, new_n19003, new_n19004, new_n19005,
    new_n19006, new_n19007, new_n19008, new_n19009, new_n19010, new_n19011,
    new_n19012, new_n19013, new_n19014, new_n19015, new_n19016, new_n19017,
    new_n19018, new_n19019, new_n19020, new_n19021, new_n19022, new_n19023,
    new_n19024, new_n19025, new_n19026, new_n19027, new_n19028, new_n19029,
    new_n19030, new_n19031, new_n19032, new_n19033, new_n19034, new_n19035,
    new_n19036, new_n19037, new_n19038, new_n19039, new_n19040, new_n19041,
    new_n19042, new_n19043, new_n19044, new_n19045, new_n19046, new_n19047,
    new_n19048, new_n19049, new_n19050, new_n19051, new_n19052, new_n19053,
    new_n19054, new_n19055, new_n19056, new_n19057, new_n19058, new_n19059,
    new_n19060, new_n19061, new_n19062, new_n19063, new_n19064, new_n19065,
    new_n19066, new_n19067, new_n19068, new_n19069, new_n19070, new_n19071,
    new_n19072, new_n19073, new_n19074, new_n19075, new_n19076, new_n19077,
    new_n19078, new_n19079, new_n19080, new_n19081, new_n19082, new_n19083,
    new_n19084, new_n19085, new_n19086, new_n19087, new_n19088, new_n19089,
    new_n19090, new_n19091, new_n19092, new_n19093, new_n19094, new_n19095,
    new_n19096, new_n19097, new_n19098, new_n19099, new_n19100, new_n19101,
    new_n19102, new_n19103, new_n19104, new_n19105, new_n19106, new_n19107,
    new_n19108, new_n19109, new_n19110, new_n19111, new_n19112, new_n19113,
    new_n19114, new_n19115, new_n19116, new_n19117, new_n19118, new_n19119,
    new_n19120, new_n19121, new_n19122, new_n19123, new_n19124, new_n19125,
    new_n19126, new_n19127, new_n19128, new_n19129, new_n19130, new_n19131,
    new_n19132, new_n19133, new_n19134, new_n19135, new_n19136, new_n19137,
    new_n19138, new_n19139, new_n19140, new_n19141, new_n19142, new_n19143,
    new_n19144, new_n19145, new_n19146, new_n19147, new_n19148, new_n19149,
    new_n19150, new_n19151, new_n19152, new_n19153, new_n19154, new_n19155,
    new_n19156, new_n19157, new_n19158, new_n19159, new_n19160, new_n19161,
    new_n19162, new_n19163, new_n19164, new_n19165, new_n19166, new_n19167,
    new_n19168, new_n19169, new_n19170, new_n19171, new_n19173, new_n19174,
    new_n19175, new_n19176, new_n19177, new_n19178, new_n19179, new_n19180,
    new_n19181, new_n19182, new_n19183, new_n19184, new_n19185, new_n19186,
    new_n19187, new_n19188, new_n19189, new_n19190, new_n19191, new_n19192,
    new_n19193, new_n19194, new_n19195, new_n19196, new_n19197, new_n19198,
    new_n19199, new_n19200, new_n19201, new_n19202, new_n19203, new_n19204,
    new_n19205, new_n19206, new_n19207, new_n19208, new_n19209, new_n19210,
    new_n19211, new_n19212, new_n19213, new_n19214, new_n19215, new_n19216,
    new_n19217, new_n19218, new_n19219, new_n19220, new_n19221, new_n19222,
    new_n19223, new_n19224, new_n19225, new_n19226, new_n19227, new_n19228,
    new_n19229, new_n19230, new_n19231, new_n19232, new_n19233, new_n19234,
    new_n19235, new_n19236, new_n19237, new_n19238, new_n19239, new_n19240,
    new_n19241, new_n19242, new_n19243, new_n19244, new_n19245, new_n19246,
    new_n19247, new_n19248, new_n19249, new_n19250, new_n19251, new_n19252,
    new_n19253, new_n19254, new_n19255, new_n19256, new_n19257, new_n19258,
    new_n19259, new_n19260, new_n19261, new_n19262, new_n19263, new_n19264,
    new_n19265, new_n19266, new_n19267, new_n19268, new_n19269, new_n19270,
    new_n19271, new_n19272, new_n19273, new_n19274, new_n19275, new_n19276,
    new_n19277, new_n19278, new_n19279, new_n19280, new_n19281, new_n19282,
    new_n19283, new_n19284, new_n19285, new_n19286, new_n19287, new_n19288,
    new_n19289, new_n19290, new_n19291, new_n19292, new_n19293, new_n19294,
    new_n19295, new_n19296, new_n19297, new_n19298, new_n19299, new_n19300,
    new_n19301, new_n19302, new_n19303, new_n19304, new_n19305, new_n19306,
    new_n19307, new_n19308, new_n19309, new_n19310, new_n19311, new_n19312,
    new_n19313, new_n19314, new_n19315, new_n19316, new_n19317, new_n19318,
    new_n19319, new_n19320, new_n19321, new_n19322, new_n19323, new_n19324,
    new_n19325, new_n19326, new_n19327, new_n19328, new_n19329, new_n19330,
    new_n19331, new_n19332, new_n19333, new_n19334, new_n19335, new_n19336,
    new_n19337, new_n19338, new_n19339, new_n19340, new_n19341, new_n19342,
    new_n19343, new_n19344, new_n19345, new_n19346, new_n19347, new_n19348,
    new_n19349, new_n19350, new_n19351, new_n19352, new_n19353, new_n19354,
    new_n19355, new_n19356, new_n19357, new_n19358, new_n19359, new_n19360,
    new_n19361, new_n19362, new_n19363, new_n19364, new_n19365, new_n19366,
    new_n19367, new_n19368, new_n19369, new_n19370, new_n19371, new_n19372,
    new_n19373, new_n19374, new_n19375, new_n19376, new_n19377, new_n19378,
    new_n19379, new_n19380, new_n19381, new_n19382, new_n19383, new_n19384,
    new_n19385, new_n19386, new_n19387, new_n19389, new_n19390, new_n19391,
    new_n19392, new_n19393, new_n19394, new_n19395, new_n19396, new_n19397,
    new_n19398, new_n19399, new_n19400, new_n19401, new_n19402, new_n19403,
    new_n19404, new_n19405, new_n19406, new_n19407, new_n19408, new_n19409,
    new_n19410, new_n19411, new_n19412, new_n19413, new_n19414, new_n19415,
    new_n19416, new_n19417, new_n19418, new_n19419, new_n19420, new_n19421,
    new_n19422, new_n19423, new_n19424, new_n19425, new_n19426, new_n19427,
    new_n19428, new_n19429, new_n19430, new_n19431, new_n19432, new_n19433,
    new_n19434, new_n19435, new_n19436, new_n19437, new_n19438, new_n19439,
    new_n19440, new_n19441, new_n19442, new_n19443, new_n19444, new_n19445,
    new_n19446, new_n19447, new_n19448, new_n19449, new_n19450, new_n19451,
    new_n19452, new_n19453, new_n19454, new_n19455, new_n19456, new_n19457,
    new_n19458, new_n19459, new_n19460, new_n19461, new_n19462, new_n19463,
    new_n19464, new_n19465, new_n19466, new_n19467, new_n19468, new_n19469,
    new_n19470, new_n19471, new_n19472, new_n19473, new_n19474, new_n19475,
    new_n19476, new_n19477, new_n19478, new_n19479, new_n19480, new_n19481,
    new_n19482, new_n19483, new_n19484, new_n19485, new_n19486, new_n19487,
    new_n19488, new_n19489, new_n19490, new_n19491, new_n19492, new_n19493,
    new_n19494, new_n19495, new_n19496, new_n19497, new_n19498, new_n19499,
    new_n19500, new_n19501, new_n19502, new_n19503, new_n19504, new_n19505,
    new_n19506, new_n19507, new_n19508, new_n19509, new_n19510, new_n19511,
    new_n19512, new_n19513, new_n19514, new_n19515, new_n19516, new_n19517,
    new_n19518, new_n19519, new_n19520, new_n19521, new_n19522, new_n19523,
    new_n19524, new_n19525, new_n19526, new_n19527, new_n19528, new_n19529,
    new_n19530, new_n19531, new_n19532, new_n19533, new_n19534, new_n19535,
    new_n19536, new_n19537, new_n19538, new_n19539, new_n19540, new_n19541,
    new_n19542, new_n19543, new_n19544, new_n19545, new_n19546, new_n19547,
    new_n19548, new_n19549, new_n19550, new_n19551, new_n19552, new_n19553,
    new_n19554, new_n19555, new_n19556, new_n19557, new_n19558, new_n19559,
    new_n19560, new_n19561, new_n19562, new_n19563, new_n19564, new_n19565,
    new_n19566, new_n19567, new_n19568, new_n19569, new_n19570, new_n19571,
    new_n19572, new_n19573, new_n19574, new_n19575, new_n19576, new_n19577,
    new_n19578, new_n19579, new_n19580, new_n19581, new_n19582, new_n19583,
    new_n19584, new_n19585, new_n19586, new_n19587, new_n19588, new_n19589,
    new_n19590, new_n19591, new_n19592, new_n19593, new_n19594, new_n19595,
    new_n19596, new_n19597, new_n19598, new_n19599, new_n19600, new_n19601,
    new_n19602, new_n19603, new_n19605, new_n19606, new_n19607, new_n19608,
    new_n19609, new_n19610, new_n19611, new_n19612, new_n19613, new_n19614,
    new_n19615, new_n19616, new_n19617, new_n19618, new_n19619, new_n19620,
    new_n19621, new_n19622, new_n19623, new_n19624, new_n19625, new_n19626,
    new_n19627, new_n19628, new_n19629, new_n19630, new_n19631, new_n19632,
    new_n19633, new_n19634, new_n19635, new_n19636, new_n19637, new_n19638,
    new_n19639, new_n19640, new_n19641, new_n19642, new_n19643, new_n19644,
    new_n19645, new_n19646, new_n19647, new_n19648, new_n19649, new_n19650,
    new_n19651, new_n19652, new_n19653, new_n19654, new_n19655, new_n19656,
    new_n19657, new_n19658, new_n19659, new_n19660, new_n19661, new_n19662,
    new_n19663, new_n19664, new_n19665, new_n19666, new_n19667, new_n19668,
    new_n19669, new_n19670, new_n19671, new_n19672, new_n19673, new_n19674,
    new_n19675, new_n19676, new_n19677, new_n19678, new_n19679, new_n19680,
    new_n19681, new_n19682, new_n19683, new_n19684, new_n19685, new_n19686,
    new_n19687, new_n19688, new_n19689, new_n19690, new_n19691, new_n19692,
    new_n19693, new_n19694, new_n19695, new_n19696, new_n19697, new_n19698,
    new_n19699, new_n19700, new_n19701, new_n19702, new_n19703, new_n19704,
    new_n19705, new_n19706, new_n19707, new_n19708, new_n19709, new_n19710,
    new_n19711, new_n19712, new_n19713, new_n19714, new_n19715, new_n19716,
    new_n19717, new_n19718, new_n19719, new_n19720, new_n19721, new_n19722,
    new_n19723, new_n19724, new_n19725, new_n19726, new_n19727, new_n19728,
    new_n19729, new_n19730, new_n19731, new_n19732, new_n19733, new_n19734,
    new_n19735, new_n19736, new_n19737, new_n19738, new_n19739, new_n19740,
    new_n19741, new_n19742, new_n19743, new_n19744, new_n19745, new_n19746,
    new_n19747, new_n19748, new_n19749, new_n19750, new_n19751, new_n19752,
    new_n19753, new_n19754, new_n19755, new_n19756, new_n19757, new_n19758,
    new_n19759, new_n19760, new_n19761, new_n19762, new_n19763, new_n19764,
    new_n19765, new_n19766, new_n19767, new_n19768, new_n19769, new_n19770,
    new_n19771, new_n19772, new_n19773, new_n19774, new_n19775, new_n19776,
    new_n19777, new_n19778, new_n19779, new_n19780, new_n19781, new_n19782,
    new_n19783, new_n19784, new_n19785, new_n19786, new_n19787, new_n19788,
    new_n19789, new_n19790, new_n19791, new_n19792, new_n19793, new_n19794,
    new_n19795, new_n19796, new_n19797, new_n19798, new_n19799, new_n19800,
    new_n19801, new_n19802, new_n19803, new_n19804, new_n19805, new_n19806,
    new_n19808, new_n19809, new_n19810, new_n19811, new_n19812, new_n19813,
    new_n19814, new_n19815, new_n19816, new_n19817, new_n19818, new_n19819,
    new_n19820, new_n19821, new_n19822, new_n19823, new_n19824, new_n19825,
    new_n19826, new_n19827, new_n19828, new_n19829, new_n19830, new_n19831,
    new_n19832, new_n19833, new_n19834, new_n19835, new_n19836, new_n19837,
    new_n19838, new_n19839, new_n19840, new_n19841, new_n19842, new_n19843,
    new_n19844, new_n19845, new_n19846, new_n19847, new_n19848, new_n19849,
    new_n19850, new_n19851, new_n19852, new_n19853, new_n19854, new_n19855,
    new_n19856, new_n19857, new_n19858, new_n19859, new_n19860, new_n19861,
    new_n19862, new_n19863, new_n19864, new_n19865, new_n19866, new_n19867,
    new_n19868, new_n19869, new_n19870, new_n19871, new_n19872, new_n19873,
    new_n19874, new_n19875, new_n19876, new_n19877, new_n19878, new_n19879,
    new_n19880, new_n19881, new_n19882, new_n19883, new_n19884, new_n19885,
    new_n19886, new_n19887, new_n19888, new_n19889, new_n19890, new_n19891,
    new_n19892, new_n19893, new_n19894, new_n19895, new_n19896, new_n19897,
    new_n19898, new_n19899, new_n19900, new_n19901, new_n19902, new_n19903,
    new_n19904, new_n19905, new_n19906, new_n19907, new_n19908, new_n19909,
    new_n19910, new_n19911, new_n19912, new_n19913, new_n19914, new_n19915,
    new_n19916, new_n19917, new_n19918, new_n19919, new_n19920, new_n19921,
    new_n19922, new_n19923, new_n19924, new_n19925, new_n19926, new_n19927,
    new_n19928, new_n19929, new_n19930, new_n19931, new_n19932, new_n19933,
    new_n19934, new_n19935, new_n19936, new_n19937, new_n19938, new_n19939,
    new_n19940, new_n19941, new_n19942, new_n19943, new_n19944, new_n19945,
    new_n19946, new_n19947, new_n19948, new_n19949, new_n19950, new_n19951,
    new_n19952, new_n19953, new_n19954, new_n19955, new_n19956, new_n19957,
    new_n19958, new_n19959, new_n19960, new_n19961, new_n19962, new_n19963,
    new_n19964, new_n19965, new_n19966, new_n19967, new_n19968, new_n19969,
    new_n19970, new_n19971, new_n19972, new_n19973, new_n19974, new_n19975,
    new_n19976, new_n19977, new_n19978, new_n19979, new_n19980, new_n19981,
    new_n19982, new_n19983, new_n19984, new_n19985, new_n19986, new_n19987,
    new_n19988, new_n19989, new_n19990, new_n19991, new_n19992, new_n19993,
    new_n19994, new_n19995, new_n19996, new_n19997, new_n19998, new_n19999,
    new_n20000, new_n20001, new_n20002, new_n20003, new_n20004, new_n20005,
    new_n20007, new_n20008, new_n20009, new_n20010, new_n20011, new_n20012,
    new_n20013, new_n20014, new_n20015, new_n20016, new_n20017, new_n20018,
    new_n20019, new_n20020, new_n20021, new_n20022, new_n20023, new_n20024,
    new_n20025, new_n20026, new_n20027, new_n20028, new_n20029, new_n20030,
    new_n20031, new_n20032, new_n20033, new_n20034, new_n20035, new_n20036,
    new_n20037, new_n20038, new_n20039, new_n20040, new_n20041, new_n20042,
    new_n20043, new_n20044, new_n20045, new_n20046, new_n20047, new_n20048,
    new_n20049, new_n20050, new_n20051, new_n20052, new_n20053, new_n20054,
    new_n20055, new_n20056, new_n20057, new_n20058, new_n20059, new_n20060,
    new_n20061, new_n20062, new_n20063, new_n20064, new_n20065, new_n20066,
    new_n20067, new_n20068, new_n20069, new_n20070, new_n20071, new_n20072,
    new_n20073, new_n20074, new_n20075, new_n20076, new_n20077, new_n20078,
    new_n20079, new_n20080, new_n20081, new_n20082, new_n20083, new_n20084,
    new_n20085, new_n20086, new_n20087, new_n20088, new_n20089, new_n20090,
    new_n20091, new_n20092, new_n20093, new_n20094, new_n20095, new_n20096,
    new_n20097, new_n20098, new_n20099, new_n20100, new_n20101, new_n20102,
    new_n20103, new_n20104, new_n20105, new_n20106, new_n20107, new_n20108,
    new_n20109, new_n20110, new_n20111, new_n20112, new_n20113, new_n20114,
    new_n20115, new_n20116, new_n20117, new_n20118, new_n20119, new_n20120,
    new_n20121, new_n20122, new_n20123, new_n20124, new_n20125, new_n20126,
    new_n20127, new_n20128, new_n20129, new_n20130, new_n20131, new_n20132,
    new_n20133, new_n20134, new_n20135, new_n20136, new_n20137, new_n20138,
    new_n20139, new_n20140, new_n20141, new_n20142, new_n20143, new_n20144,
    new_n20145, new_n20146, new_n20147, new_n20148, new_n20149, new_n20150,
    new_n20151, new_n20152, new_n20153, new_n20154, new_n20155, new_n20156,
    new_n20157, new_n20158, new_n20159, new_n20160, new_n20161, new_n20162,
    new_n20163, new_n20164, new_n20165, new_n20166, new_n20167, new_n20168,
    new_n20169, new_n20170, new_n20171, new_n20172, new_n20173, new_n20174,
    new_n20175, new_n20176, new_n20177, new_n20178, new_n20179, new_n20180,
    new_n20181, new_n20182, new_n20183, new_n20184, new_n20185, new_n20186,
    new_n20187, new_n20188, new_n20189, new_n20190, new_n20191, new_n20192,
    new_n20193, new_n20194, new_n20195, new_n20196, new_n20197, new_n20198,
    new_n20199, new_n20200, new_n20202, new_n20203, new_n20204, new_n20205,
    new_n20206, new_n20207, new_n20208, new_n20209, new_n20210, new_n20211,
    new_n20212, new_n20213, new_n20214, new_n20215, new_n20216, new_n20217,
    new_n20218, new_n20219, new_n20220, new_n20221, new_n20222, new_n20223,
    new_n20224, new_n20225, new_n20226, new_n20227, new_n20228, new_n20229,
    new_n20230, new_n20231, new_n20232, new_n20233, new_n20234, new_n20235,
    new_n20236, new_n20237, new_n20238, new_n20239, new_n20240, new_n20241,
    new_n20242, new_n20243, new_n20244, new_n20245, new_n20246, new_n20247,
    new_n20248, new_n20249, new_n20250, new_n20251, new_n20252, new_n20253,
    new_n20254, new_n20255, new_n20256, new_n20257, new_n20258, new_n20259,
    new_n20260, new_n20261, new_n20262, new_n20263, new_n20264, new_n20265,
    new_n20266, new_n20267, new_n20268, new_n20269, new_n20270, new_n20271,
    new_n20272, new_n20273, new_n20274, new_n20275, new_n20276, new_n20277,
    new_n20278, new_n20279, new_n20280, new_n20281, new_n20282, new_n20283,
    new_n20284, new_n20285, new_n20286, new_n20287, new_n20288, new_n20289,
    new_n20290, new_n20291, new_n20292, new_n20293, new_n20294, new_n20295,
    new_n20296, new_n20297, new_n20298, new_n20299, new_n20300, new_n20301,
    new_n20302, new_n20303, new_n20304, new_n20305, new_n20306, new_n20307,
    new_n20308, new_n20309, new_n20310, new_n20311, new_n20312, new_n20313,
    new_n20314, new_n20315, new_n20316, new_n20317, new_n20318, new_n20319,
    new_n20320, new_n20321, new_n20322, new_n20323, new_n20324, new_n20325,
    new_n20326, new_n20327, new_n20328, new_n20329, new_n20330, new_n20331,
    new_n20332, new_n20333, new_n20334, new_n20335, new_n20336, new_n20337,
    new_n20338, new_n20339, new_n20340, new_n20341, new_n20342, new_n20343,
    new_n20344, new_n20345, new_n20346, new_n20347, new_n20348, new_n20349,
    new_n20350, new_n20351, new_n20352, new_n20353, new_n20354, new_n20355,
    new_n20356, new_n20357, new_n20358, new_n20359, new_n20360, new_n20361,
    new_n20362, new_n20363, new_n20364, new_n20365, new_n20366, new_n20367,
    new_n20368, new_n20369, new_n20370, new_n20371, new_n20372, new_n20373,
    new_n20374, new_n20375, new_n20376, new_n20377, new_n20378, new_n20379,
    new_n20380, new_n20381, new_n20382, new_n20383, new_n20384, new_n20385,
    new_n20386, new_n20387, new_n20388, new_n20389, new_n20391, new_n20392,
    new_n20393, new_n20394, new_n20395, new_n20396, new_n20397, new_n20398,
    new_n20399, new_n20400, new_n20401, new_n20402, new_n20403, new_n20404,
    new_n20405, new_n20406, new_n20407, new_n20408, new_n20409, new_n20410,
    new_n20411, new_n20412, new_n20413, new_n20414, new_n20415, new_n20416,
    new_n20417, new_n20418, new_n20419, new_n20420, new_n20421, new_n20422,
    new_n20423, new_n20424, new_n20425, new_n20426, new_n20427, new_n20428,
    new_n20429, new_n20430, new_n20431, new_n20432, new_n20433, new_n20434,
    new_n20435, new_n20436, new_n20437, new_n20438, new_n20439, new_n20440,
    new_n20441, new_n20442, new_n20443, new_n20444, new_n20445, new_n20446,
    new_n20447, new_n20448, new_n20449, new_n20450, new_n20451, new_n20452,
    new_n20453, new_n20454, new_n20455, new_n20456, new_n20457, new_n20458,
    new_n20459, new_n20460, new_n20461, new_n20462, new_n20463, new_n20464,
    new_n20465, new_n20466, new_n20467, new_n20468, new_n20469, new_n20470,
    new_n20471, new_n20472, new_n20473, new_n20474, new_n20475, new_n20476,
    new_n20477, new_n20478, new_n20479, new_n20480, new_n20481, new_n20482,
    new_n20483, new_n20484, new_n20485, new_n20486, new_n20487, new_n20488,
    new_n20489, new_n20490, new_n20491, new_n20492, new_n20493, new_n20494,
    new_n20495, new_n20496, new_n20497, new_n20498, new_n20499, new_n20500,
    new_n20501, new_n20502, new_n20503, new_n20504, new_n20505, new_n20506,
    new_n20507, new_n20508, new_n20509, new_n20510, new_n20511, new_n20512,
    new_n20513, new_n20514, new_n20515, new_n20516, new_n20517, new_n20518,
    new_n20519, new_n20520, new_n20521, new_n20522, new_n20523, new_n20524,
    new_n20525, new_n20526, new_n20527, new_n20528, new_n20529, new_n20530,
    new_n20531, new_n20532, new_n20533, new_n20534, new_n20535, new_n20536,
    new_n20537, new_n20538, new_n20539, new_n20540, new_n20541, new_n20542,
    new_n20543, new_n20544, new_n20545, new_n20546, new_n20547, new_n20548,
    new_n20549, new_n20550, new_n20551, new_n20552, new_n20553, new_n20554,
    new_n20555, new_n20556, new_n20557, new_n20558, new_n20559, new_n20560,
    new_n20561, new_n20562, new_n20563, new_n20564, new_n20565, new_n20566,
    new_n20567, new_n20568, new_n20569, new_n20570, new_n20571, new_n20572,
    new_n20573, new_n20574, new_n20575, new_n20576, new_n20578, new_n20579,
    new_n20580, new_n20581, new_n20582, new_n20583, new_n20584, new_n20585,
    new_n20586, new_n20587, new_n20588, new_n20589, new_n20590, new_n20591,
    new_n20592, new_n20593, new_n20594, new_n20595, new_n20596, new_n20597,
    new_n20598, new_n20599, new_n20600, new_n20601, new_n20602, new_n20603,
    new_n20604, new_n20605, new_n20606, new_n20607, new_n20608, new_n20609,
    new_n20610, new_n20611, new_n20612, new_n20613, new_n20614, new_n20615,
    new_n20616, new_n20617, new_n20618, new_n20619, new_n20620, new_n20621,
    new_n20622, new_n20623, new_n20624, new_n20625, new_n20626, new_n20627,
    new_n20628, new_n20629, new_n20630, new_n20631, new_n20632, new_n20633,
    new_n20634, new_n20635, new_n20636, new_n20637, new_n20638, new_n20639,
    new_n20640, new_n20641, new_n20642, new_n20643, new_n20644, new_n20645,
    new_n20646, new_n20647, new_n20648, new_n20649, new_n20650, new_n20651,
    new_n20652, new_n20653, new_n20654, new_n20655, new_n20656, new_n20657,
    new_n20658, new_n20659, new_n20660, new_n20661, new_n20662, new_n20663,
    new_n20664, new_n20665, new_n20666, new_n20667, new_n20668, new_n20669,
    new_n20670, new_n20671, new_n20672, new_n20673, new_n20674, new_n20675,
    new_n20676, new_n20677, new_n20678, new_n20679, new_n20680, new_n20681,
    new_n20682, new_n20683, new_n20684, new_n20685, new_n20686, new_n20687,
    new_n20688, new_n20689, new_n20690, new_n20691, new_n20692, new_n20693,
    new_n20694, new_n20695, new_n20696, new_n20697, new_n20698, new_n20699,
    new_n20700, new_n20701, new_n20702, new_n20703, new_n20704, new_n20705,
    new_n20706, new_n20707, new_n20708, new_n20709, new_n20710, new_n20711,
    new_n20712, new_n20713, new_n20714, new_n20715, new_n20716, new_n20717,
    new_n20718, new_n20719, new_n20720, new_n20721, new_n20722, new_n20723,
    new_n20724, new_n20725, new_n20726, new_n20727, new_n20728, new_n20729,
    new_n20730, new_n20731, new_n20732, new_n20733, new_n20734, new_n20735,
    new_n20736, new_n20737, new_n20738, new_n20739, new_n20740, new_n20741,
    new_n20742, new_n20743, new_n20744, new_n20745, new_n20746, new_n20747,
    new_n20748, new_n20749, new_n20750, new_n20751, new_n20752, new_n20753,
    new_n20755, new_n20756, new_n20757, new_n20758, new_n20759, new_n20760,
    new_n20761, new_n20762, new_n20763, new_n20764, new_n20765, new_n20766,
    new_n20767, new_n20768, new_n20769, new_n20770, new_n20771, new_n20772,
    new_n20773, new_n20774, new_n20775, new_n20776, new_n20777, new_n20778,
    new_n20779, new_n20780, new_n20781, new_n20782, new_n20783, new_n20784,
    new_n20785, new_n20786, new_n20787, new_n20788, new_n20789, new_n20790,
    new_n20791, new_n20792, new_n20793, new_n20794, new_n20795, new_n20796,
    new_n20797, new_n20798, new_n20799, new_n20800, new_n20801, new_n20802,
    new_n20803, new_n20804, new_n20805, new_n20806, new_n20807, new_n20808,
    new_n20809, new_n20810, new_n20811, new_n20812, new_n20813, new_n20814,
    new_n20815, new_n20816, new_n20817, new_n20818, new_n20819, new_n20820,
    new_n20821, new_n20822, new_n20823, new_n20824, new_n20825, new_n20826,
    new_n20827, new_n20828, new_n20829, new_n20830, new_n20831, new_n20832,
    new_n20833, new_n20834, new_n20835, new_n20836, new_n20837, new_n20838,
    new_n20839, new_n20840, new_n20841, new_n20842, new_n20843, new_n20844,
    new_n20845, new_n20846, new_n20847, new_n20848, new_n20849, new_n20850,
    new_n20851, new_n20852, new_n20853, new_n20854, new_n20855, new_n20856,
    new_n20857, new_n20858, new_n20859, new_n20860, new_n20861, new_n20862,
    new_n20863, new_n20864, new_n20865, new_n20866, new_n20867, new_n20868,
    new_n20869, new_n20870, new_n20871, new_n20872, new_n20873, new_n20874,
    new_n20875, new_n20876, new_n20877, new_n20878, new_n20879, new_n20880,
    new_n20881, new_n20882, new_n20883, new_n20884, new_n20885, new_n20886,
    new_n20887, new_n20888, new_n20889, new_n20890, new_n20891, new_n20892,
    new_n20893, new_n20894, new_n20895, new_n20896, new_n20897, new_n20898,
    new_n20899, new_n20900, new_n20901, new_n20902, new_n20903, new_n20904,
    new_n20905, new_n20906, new_n20907, new_n20908, new_n20909, new_n20910,
    new_n20911, new_n20912, new_n20913, new_n20914, new_n20915, new_n20916,
    new_n20917, new_n20918, new_n20919, new_n20920, new_n20922, new_n20923,
    new_n20924, new_n20925, new_n20926, new_n20927, new_n20928, new_n20929,
    new_n20930, new_n20931, new_n20932, new_n20933, new_n20934, new_n20935,
    new_n20936, new_n20937, new_n20938, new_n20939, new_n20940, new_n20941,
    new_n20942, new_n20943, new_n20944, new_n20945, new_n20946, new_n20947,
    new_n20948, new_n20949, new_n20950, new_n20951, new_n20952, new_n20953,
    new_n20954, new_n20955, new_n20956, new_n20957, new_n20958, new_n20959,
    new_n20960, new_n20961, new_n20962, new_n20963, new_n20964, new_n20965,
    new_n20966, new_n20967, new_n20968, new_n20969, new_n20970, new_n20971,
    new_n20972, new_n20973, new_n20974, new_n20975, new_n20976, new_n20977,
    new_n20978, new_n20979, new_n20980, new_n20981, new_n20982, new_n20983,
    new_n20984, new_n20985, new_n20986, new_n20987, new_n20988, new_n20989,
    new_n20990, new_n20991, new_n20992, new_n20993, new_n20994, new_n20995,
    new_n20996, new_n20997, new_n20998, new_n20999, new_n21000, new_n21001,
    new_n21002, new_n21003, new_n21004, new_n21005, new_n21006, new_n21007,
    new_n21008, new_n21009, new_n21010, new_n21011, new_n21012, new_n21013,
    new_n21014, new_n21015, new_n21016, new_n21017, new_n21018, new_n21019,
    new_n21020, new_n21021, new_n21022, new_n21023, new_n21024, new_n21025,
    new_n21026, new_n21027, new_n21028, new_n21029, new_n21030, new_n21031,
    new_n21032, new_n21033, new_n21034, new_n21035, new_n21036, new_n21037,
    new_n21038, new_n21039, new_n21040, new_n21041, new_n21042, new_n21043,
    new_n21044, new_n21045, new_n21046, new_n21047, new_n21048, new_n21049,
    new_n21050, new_n21051, new_n21052, new_n21053, new_n21054, new_n21055,
    new_n21056, new_n21057, new_n21058, new_n21059, new_n21060, new_n21061,
    new_n21062, new_n21063, new_n21064, new_n21065, new_n21066, new_n21067,
    new_n21068, new_n21069, new_n21070, new_n21071, new_n21072, new_n21073,
    new_n21074, new_n21075, new_n21076, new_n21077, new_n21078, new_n21079,
    new_n21080, new_n21081, new_n21082, new_n21083, new_n21085, new_n21086,
    new_n21087, new_n21088, new_n21089, new_n21090, new_n21091, new_n21092,
    new_n21093, new_n21094, new_n21095, new_n21096, new_n21097, new_n21098,
    new_n21099, new_n21100, new_n21101, new_n21102, new_n21103, new_n21104,
    new_n21105, new_n21106, new_n21107, new_n21108, new_n21109, new_n21110,
    new_n21111, new_n21112, new_n21113, new_n21114, new_n21115, new_n21116,
    new_n21117, new_n21118, new_n21119, new_n21120, new_n21121, new_n21122,
    new_n21123, new_n21124, new_n21125, new_n21126, new_n21127, new_n21128,
    new_n21129, new_n21130, new_n21131, new_n21132, new_n21133, new_n21134,
    new_n21135, new_n21136, new_n21137, new_n21138, new_n21139, new_n21140,
    new_n21141, new_n21142, new_n21143, new_n21144, new_n21145, new_n21146,
    new_n21147, new_n21148, new_n21149, new_n21150, new_n21151, new_n21152,
    new_n21153, new_n21154, new_n21155, new_n21156, new_n21157, new_n21158,
    new_n21159, new_n21160, new_n21161, new_n21162, new_n21163, new_n21164,
    new_n21165, new_n21166, new_n21167, new_n21168, new_n21169, new_n21170,
    new_n21171, new_n21172, new_n21173, new_n21174, new_n21175, new_n21176,
    new_n21177, new_n21178, new_n21179, new_n21180, new_n21181, new_n21182,
    new_n21183, new_n21184, new_n21185, new_n21186, new_n21187, new_n21188,
    new_n21189, new_n21190, new_n21191, new_n21192, new_n21193, new_n21194,
    new_n21195, new_n21196, new_n21197, new_n21198, new_n21199, new_n21200,
    new_n21201, new_n21202, new_n21203, new_n21204, new_n21205, new_n21206,
    new_n21207, new_n21208, new_n21209, new_n21210, new_n21211, new_n21212,
    new_n21213, new_n21214, new_n21215, new_n21216, new_n21217, new_n21218,
    new_n21219, new_n21220, new_n21221, new_n21222, new_n21223, new_n21224,
    new_n21225, new_n21226, new_n21227, new_n21228, new_n21229, new_n21230,
    new_n21231, new_n21232, new_n21233, new_n21234, new_n21235, new_n21236,
    new_n21237, new_n21238, new_n21240, new_n21241, new_n21242, new_n21243,
    new_n21244, new_n21245, new_n21246, new_n21247, new_n21248, new_n21249,
    new_n21250, new_n21251, new_n21252, new_n21253, new_n21254, new_n21255,
    new_n21256, new_n21257, new_n21258, new_n21259, new_n21260, new_n21261,
    new_n21262, new_n21263, new_n21264, new_n21265, new_n21266, new_n21267,
    new_n21268, new_n21269, new_n21270, new_n21271, new_n21272, new_n21273,
    new_n21274, new_n21275, new_n21276, new_n21277, new_n21278, new_n21279,
    new_n21280, new_n21281, new_n21282, new_n21283, new_n21284, new_n21285,
    new_n21286, new_n21287, new_n21288, new_n21289, new_n21290, new_n21291,
    new_n21292, new_n21293, new_n21294, new_n21295, new_n21296, new_n21297,
    new_n21298, new_n21299, new_n21300, new_n21301, new_n21302, new_n21303,
    new_n21304, new_n21305, new_n21306, new_n21307, new_n21308, new_n21309,
    new_n21310, new_n21311, new_n21312, new_n21313, new_n21314, new_n21315,
    new_n21316, new_n21317, new_n21318, new_n21319, new_n21320, new_n21321,
    new_n21322, new_n21323, new_n21324, new_n21325, new_n21326, new_n21327,
    new_n21328, new_n21329, new_n21330, new_n21331, new_n21332, new_n21333,
    new_n21334, new_n21335, new_n21336, new_n21337, new_n21338, new_n21339,
    new_n21340, new_n21341, new_n21342, new_n21343, new_n21344, new_n21345,
    new_n21346, new_n21347, new_n21348, new_n21349, new_n21350, new_n21351,
    new_n21352, new_n21353, new_n21354, new_n21355, new_n21356, new_n21357,
    new_n21358, new_n21359, new_n21360, new_n21361, new_n21362, new_n21363,
    new_n21364, new_n21365, new_n21366, new_n21367, new_n21368, new_n21369,
    new_n21370, new_n21371, new_n21372, new_n21373, new_n21374, new_n21375,
    new_n21376, new_n21377, new_n21378, new_n21379, new_n21380, new_n21381,
    new_n21382, new_n21383, new_n21384, new_n21385, new_n21386, new_n21387,
    new_n21388, new_n21389, new_n21390, new_n21392, new_n21393, new_n21394,
    new_n21395, new_n21396, new_n21397, new_n21398, new_n21399, new_n21400,
    new_n21401, new_n21402, new_n21403, new_n21404, new_n21405, new_n21406,
    new_n21407, new_n21408, new_n21409, new_n21410, new_n21411, new_n21412,
    new_n21413, new_n21414, new_n21415, new_n21416, new_n21417, new_n21418,
    new_n21419, new_n21420, new_n21421, new_n21422, new_n21423, new_n21424,
    new_n21425, new_n21426, new_n21427, new_n21428, new_n21429, new_n21430,
    new_n21431, new_n21432, new_n21433, new_n21434, new_n21435, new_n21436,
    new_n21437, new_n21438, new_n21439, new_n21440, new_n21441, new_n21442,
    new_n21443, new_n21444, new_n21445, new_n21446, new_n21447, new_n21448,
    new_n21449, new_n21450, new_n21451, new_n21452, new_n21453, new_n21454,
    new_n21455, new_n21456, new_n21457, new_n21458, new_n21459, new_n21460,
    new_n21461, new_n21462, new_n21463, new_n21464, new_n21465, new_n21466,
    new_n21467, new_n21468, new_n21469, new_n21470, new_n21471, new_n21472,
    new_n21473, new_n21474, new_n21475, new_n21476, new_n21477, new_n21478,
    new_n21479, new_n21480, new_n21481, new_n21482, new_n21483, new_n21484,
    new_n21485, new_n21486, new_n21487, new_n21488, new_n21489, new_n21490,
    new_n21491, new_n21492, new_n21493, new_n21494, new_n21495, new_n21496,
    new_n21497, new_n21498, new_n21499, new_n21500, new_n21501, new_n21502,
    new_n21503, new_n21504, new_n21505, new_n21506, new_n21507, new_n21508,
    new_n21509, new_n21510, new_n21511, new_n21512, new_n21513, new_n21514,
    new_n21515, new_n21516, new_n21517, new_n21518, new_n21519, new_n21520,
    new_n21521, new_n21522, new_n21523, new_n21524, new_n21525, new_n21526,
    new_n21527, new_n21528, new_n21529, new_n21530, new_n21531, new_n21532,
    new_n21533, new_n21534, new_n21535, new_n21536, new_n21537, new_n21538,
    new_n21540, new_n21541, new_n21542, new_n21543, new_n21544, new_n21545,
    new_n21546, new_n21547, new_n21548, new_n21549, new_n21550, new_n21551,
    new_n21552, new_n21553, new_n21554, new_n21555, new_n21556, new_n21557,
    new_n21558, new_n21559, new_n21560, new_n21561, new_n21562, new_n21563,
    new_n21564, new_n21565, new_n21566, new_n21567, new_n21568, new_n21569,
    new_n21570, new_n21571, new_n21572, new_n21573, new_n21574, new_n21575,
    new_n21576, new_n21577, new_n21578, new_n21579, new_n21580, new_n21581,
    new_n21582, new_n21583, new_n21584, new_n21585, new_n21586, new_n21587,
    new_n21588, new_n21589, new_n21590, new_n21591, new_n21592, new_n21593,
    new_n21594, new_n21595, new_n21596, new_n21597, new_n21598, new_n21599,
    new_n21600, new_n21601, new_n21602, new_n21603, new_n21604, new_n21605,
    new_n21606, new_n21607, new_n21608, new_n21609, new_n21610, new_n21611,
    new_n21612, new_n21613, new_n21614, new_n21615, new_n21616, new_n21617,
    new_n21618, new_n21619, new_n21620, new_n21621, new_n21622, new_n21623,
    new_n21624, new_n21625, new_n21626, new_n21627, new_n21628, new_n21629,
    new_n21630, new_n21631, new_n21632, new_n21633, new_n21634, new_n21635,
    new_n21636, new_n21637, new_n21638, new_n21639, new_n21640, new_n21641,
    new_n21642, new_n21643, new_n21644, new_n21645, new_n21646, new_n21647,
    new_n21648, new_n21649, new_n21650, new_n21651, new_n21652, new_n21653,
    new_n21654, new_n21655, new_n21656, new_n21657, new_n21658, new_n21659,
    new_n21660, new_n21661, new_n21662, new_n21663, new_n21664, new_n21665,
    new_n21666, new_n21667, new_n21668, new_n21669, new_n21670, new_n21671,
    new_n21672, new_n21673, new_n21674, new_n21675, new_n21676, new_n21677,
    new_n21678, new_n21679, new_n21680, new_n21681, new_n21682, new_n21684,
    new_n21685, new_n21686, new_n21687, new_n21688, new_n21689, new_n21690,
    new_n21691, new_n21692, new_n21693, new_n21694, new_n21695, new_n21696,
    new_n21697, new_n21698, new_n21699, new_n21700, new_n21701, new_n21702,
    new_n21703, new_n21704, new_n21705, new_n21706, new_n21707, new_n21708,
    new_n21709, new_n21710, new_n21711, new_n21712, new_n21713, new_n21714,
    new_n21715, new_n21716, new_n21717, new_n21718, new_n21719, new_n21720,
    new_n21721, new_n21722, new_n21723, new_n21724, new_n21725, new_n21726,
    new_n21727, new_n21728, new_n21729, new_n21730, new_n21731, new_n21732,
    new_n21733, new_n21734, new_n21735, new_n21736, new_n21737, new_n21738,
    new_n21739, new_n21740, new_n21741, new_n21742, new_n21743, new_n21744,
    new_n21745, new_n21746, new_n21747, new_n21748, new_n21749, new_n21750,
    new_n21751, new_n21752, new_n21753, new_n21754, new_n21755, new_n21756,
    new_n21757, new_n21758, new_n21759, new_n21760, new_n21761, new_n21762,
    new_n21763, new_n21764, new_n21765, new_n21766, new_n21767, new_n21768,
    new_n21769, new_n21770, new_n21771, new_n21772, new_n21773, new_n21774,
    new_n21775, new_n21776, new_n21777, new_n21778, new_n21779, new_n21780,
    new_n21781, new_n21782, new_n21783, new_n21784, new_n21785, new_n21786,
    new_n21787, new_n21788, new_n21789, new_n21790, new_n21791, new_n21792,
    new_n21793, new_n21794, new_n21795, new_n21796, new_n21797, new_n21798,
    new_n21799, new_n21800, new_n21801, new_n21802, new_n21803, new_n21804,
    new_n21805, new_n21806, new_n21807, new_n21808, new_n21809, new_n21810,
    new_n21811, new_n21812, new_n21813, new_n21814, new_n21815, new_n21816,
    new_n21817, new_n21818, new_n21819, new_n21821, new_n21822, new_n21823,
    new_n21824, new_n21825, new_n21826, new_n21827, new_n21828, new_n21829,
    new_n21830, new_n21831, new_n21832, new_n21833, new_n21834, new_n21835,
    new_n21836, new_n21837, new_n21838, new_n21839, new_n21840, new_n21841,
    new_n21842, new_n21843, new_n21844, new_n21845, new_n21846, new_n21847,
    new_n21848, new_n21849, new_n21850, new_n21851, new_n21852, new_n21853,
    new_n21854, new_n21855, new_n21856, new_n21857, new_n21858, new_n21859,
    new_n21860, new_n21861, new_n21862, new_n21863, new_n21864, new_n21865,
    new_n21866, new_n21867, new_n21868, new_n21869, new_n21870, new_n21871,
    new_n21872, new_n21873, new_n21874, new_n21875, new_n21876, new_n21877,
    new_n21878, new_n21879, new_n21880, new_n21881, new_n21882, new_n21883,
    new_n21884, new_n21885, new_n21886, new_n21887, new_n21888, new_n21889,
    new_n21890, new_n21891, new_n21892, new_n21893, new_n21894, new_n21895,
    new_n21896, new_n21897, new_n21898, new_n21899, new_n21900, new_n21901,
    new_n21902, new_n21903, new_n21904, new_n21905, new_n21906, new_n21907,
    new_n21908, new_n21909, new_n21910, new_n21911, new_n21912, new_n21913,
    new_n21914, new_n21915, new_n21916, new_n21917, new_n21918, new_n21919,
    new_n21920, new_n21921, new_n21922, new_n21923, new_n21924, new_n21925,
    new_n21926, new_n21927, new_n21928, new_n21929, new_n21930, new_n21931,
    new_n21932, new_n21933, new_n21934, new_n21935, new_n21936, new_n21937,
    new_n21938, new_n21939, new_n21940, new_n21941, new_n21942, new_n21943,
    new_n21944, new_n21945, new_n21946, new_n21947, new_n21948, new_n21949,
    new_n21950, new_n21951, new_n21953, new_n21954, new_n21955, new_n21956,
    new_n21957, new_n21958, new_n21959, new_n21960, new_n21961, new_n21962,
    new_n21963, new_n21964, new_n21965, new_n21966, new_n21967, new_n21968,
    new_n21969, new_n21970, new_n21971, new_n21972, new_n21973, new_n21974,
    new_n21975, new_n21976, new_n21977, new_n21978, new_n21979, new_n21980,
    new_n21981, new_n21982, new_n21983, new_n21984, new_n21985, new_n21986,
    new_n21987, new_n21988, new_n21989, new_n21990, new_n21991, new_n21992,
    new_n21993, new_n21994, new_n21995, new_n21996, new_n21997, new_n21998,
    new_n21999, new_n22000, new_n22001, new_n22002, new_n22003, new_n22004,
    new_n22005, new_n22006, new_n22007, new_n22008, new_n22009, new_n22010,
    new_n22011, new_n22012, new_n22013, new_n22014, new_n22015, new_n22016,
    new_n22017, new_n22018, new_n22019, new_n22020, new_n22021, new_n22022,
    new_n22023, new_n22024, new_n22025, new_n22026, new_n22027, new_n22028,
    new_n22029, new_n22030, new_n22031, new_n22032, new_n22033, new_n22034,
    new_n22035, new_n22036, new_n22037, new_n22038, new_n22039, new_n22040,
    new_n22041, new_n22042, new_n22043, new_n22044, new_n22045, new_n22046,
    new_n22047, new_n22048, new_n22049, new_n22050, new_n22051, new_n22052,
    new_n22053, new_n22054, new_n22055, new_n22056, new_n22057, new_n22058,
    new_n22059, new_n22060, new_n22061, new_n22062, new_n22063, new_n22064,
    new_n22065, new_n22066, new_n22067, new_n22068, new_n22069, new_n22070,
    new_n22071, new_n22072, new_n22074, new_n22075, new_n22076, new_n22077,
    new_n22078, new_n22079, new_n22080, new_n22081, new_n22082, new_n22083,
    new_n22084, new_n22085, new_n22086, new_n22087, new_n22088, new_n22089,
    new_n22090, new_n22091, new_n22092, new_n22093, new_n22094, new_n22095,
    new_n22096, new_n22097, new_n22098, new_n22099, new_n22100, new_n22101,
    new_n22102, new_n22103, new_n22104, new_n22105, new_n22106, new_n22107,
    new_n22108, new_n22109, new_n22110, new_n22111, new_n22112, new_n22113,
    new_n22114, new_n22115, new_n22116, new_n22117, new_n22118, new_n22119,
    new_n22120, new_n22121, new_n22122, new_n22123, new_n22124, new_n22125,
    new_n22126, new_n22127, new_n22128, new_n22129, new_n22130, new_n22131,
    new_n22132, new_n22133, new_n22134, new_n22135, new_n22136, new_n22137,
    new_n22138, new_n22139, new_n22140, new_n22141, new_n22142, new_n22143,
    new_n22144, new_n22145, new_n22146, new_n22147, new_n22148, new_n22149,
    new_n22150, new_n22151, new_n22152, new_n22153, new_n22154, new_n22155,
    new_n22156, new_n22157, new_n22158, new_n22159, new_n22160, new_n22161,
    new_n22162, new_n22163, new_n22164, new_n22165, new_n22166, new_n22167,
    new_n22168, new_n22169, new_n22170, new_n22171, new_n22172, new_n22173,
    new_n22174, new_n22175, new_n22176, new_n22177, new_n22178, new_n22179,
    new_n22180, new_n22181, new_n22182, new_n22183, new_n22184, new_n22185,
    new_n22186, new_n22187, new_n22188, new_n22189, new_n22190, new_n22192,
    new_n22193, new_n22194, new_n22195, new_n22196, new_n22197, new_n22198,
    new_n22199, new_n22200, new_n22201, new_n22202, new_n22203, new_n22204,
    new_n22205, new_n22206, new_n22207, new_n22208, new_n22209, new_n22210,
    new_n22211, new_n22212, new_n22213, new_n22214, new_n22215, new_n22216,
    new_n22217, new_n22218, new_n22219, new_n22220, new_n22221, new_n22222,
    new_n22223, new_n22224, new_n22225, new_n22226, new_n22227, new_n22228,
    new_n22229, new_n22230, new_n22231, new_n22232, new_n22233, new_n22234,
    new_n22235, new_n22236, new_n22237, new_n22238, new_n22239, new_n22240,
    new_n22241, new_n22242, new_n22243, new_n22244, new_n22245, new_n22246,
    new_n22247, new_n22248, new_n22249, new_n22250, new_n22251, new_n22252,
    new_n22253, new_n22254, new_n22255, new_n22256, new_n22257, new_n22258,
    new_n22259, new_n22260, new_n22261, new_n22262, new_n22263, new_n22264,
    new_n22265, new_n22266, new_n22267, new_n22268, new_n22269, new_n22270,
    new_n22271, new_n22272, new_n22273, new_n22274, new_n22275, new_n22276,
    new_n22277, new_n22278, new_n22279, new_n22280, new_n22281, new_n22282,
    new_n22283, new_n22284, new_n22285, new_n22286, new_n22287, new_n22288,
    new_n22289, new_n22290, new_n22291, new_n22292, new_n22293, new_n22294,
    new_n22295, new_n22296, new_n22297, new_n22298, new_n22299, new_n22300,
    new_n22301, new_n22302, new_n22303, new_n22304, new_n22306, new_n22307,
    new_n22308, new_n22309, new_n22310, new_n22311, new_n22312, new_n22313,
    new_n22314, new_n22315, new_n22316, new_n22317, new_n22318, new_n22319,
    new_n22320, new_n22321, new_n22322, new_n22323, new_n22324, new_n22325,
    new_n22326, new_n22327, new_n22328, new_n22329, new_n22330, new_n22331,
    new_n22332, new_n22333, new_n22334, new_n22335, new_n22336, new_n22337,
    new_n22338, new_n22339, new_n22340, new_n22341, new_n22342, new_n22343,
    new_n22344, new_n22345, new_n22346, new_n22347, new_n22348, new_n22349,
    new_n22350, new_n22351, new_n22352, new_n22353, new_n22354, new_n22355,
    new_n22356, new_n22357, new_n22358, new_n22359, new_n22360, new_n22361,
    new_n22362, new_n22363, new_n22364, new_n22365, new_n22366, new_n22367,
    new_n22368, new_n22369, new_n22370, new_n22371, new_n22372, new_n22373,
    new_n22374, new_n22375, new_n22376, new_n22377, new_n22378, new_n22379,
    new_n22380, new_n22381, new_n22382, new_n22383, new_n22384, new_n22385,
    new_n22386, new_n22387, new_n22388, new_n22389, new_n22390, new_n22391,
    new_n22392, new_n22393, new_n22394, new_n22395, new_n22396, new_n22397,
    new_n22398, new_n22399, new_n22400, new_n22401, new_n22402, new_n22403,
    new_n22404, new_n22405, new_n22406, new_n22407, new_n22408, new_n22409,
    new_n22410, new_n22411, new_n22412, new_n22414, new_n22415, new_n22416,
    new_n22417, new_n22418, new_n22419, new_n22420, new_n22421, new_n22422,
    new_n22423, new_n22424, new_n22425, new_n22426, new_n22427, new_n22428,
    new_n22429, new_n22430, new_n22431, new_n22432, new_n22433, new_n22434,
    new_n22435, new_n22436, new_n22437, new_n22438, new_n22439, new_n22440,
    new_n22441, new_n22442, new_n22443, new_n22444, new_n22445, new_n22446,
    new_n22447, new_n22448, new_n22449, new_n22450, new_n22451, new_n22452,
    new_n22453, new_n22454, new_n22455, new_n22456, new_n22457, new_n22458,
    new_n22459, new_n22460, new_n22461, new_n22462, new_n22463, new_n22464,
    new_n22465, new_n22466, new_n22467, new_n22468, new_n22469, new_n22470,
    new_n22471, new_n22472, new_n22473, new_n22474, new_n22475, new_n22476,
    new_n22477, new_n22478, new_n22479, new_n22480, new_n22481, new_n22482,
    new_n22483, new_n22484, new_n22485, new_n22486, new_n22487, new_n22488,
    new_n22489, new_n22490, new_n22491, new_n22492, new_n22493, new_n22494,
    new_n22495, new_n22496, new_n22497, new_n22498, new_n22499, new_n22500,
    new_n22501, new_n22502, new_n22503, new_n22504, new_n22505, new_n22506,
    new_n22507, new_n22508, new_n22509, new_n22510, new_n22511, new_n22512,
    new_n22513, new_n22515, new_n22516, new_n22517, new_n22518, new_n22519,
    new_n22520, new_n22521, new_n22522, new_n22523, new_n22524, new_n22525,
    new_n22526, new_n22527, new_n22528, new_n22529, new_n22530, new_n22531,
    new_n22532, new_n22533, new_n22534, new_n22535, new_n22536, new_n22537,
    new_n22538, new_n22539, new_n22540, new_n22541, new_n22542, new_n22543,
    new_n22544, new_n22545, new_n22546, new_n22547, new_n22548, new_n22549,
    new_n22550, new_n22551, new_n22552, new_n22553, new_n22554, new_n22555,
    new_n22556, new_n22557, new_n22558, new_n22559, new_n22560, new_n22561,
    new_n22562, new_n22563, new_n22564, new_n22565, new_n22566, new_n22567,
    new_n22568, new_n22569, new_n22570, new_n22571, new_n22572, new_n22573,
    new_n22574, new_n22575, new_n22576, new_n22577, new_n22578, new_n22579,
    new_n22580, new_n22581, new_n22582, new_n22583, new_n22584, new_n22585,
    new_n22586, new_n22587, new_n22588, new_n22589, new_n22590, new_n22591,
    new_n22592, new_n22593, new_n22594, new_n22595, new_n22596, new_n22597,
    new_n22598, new_n22599, new_n22600, new_n22601, new_n22602, new_n22603,
    new_n22604, new_n22605, new_n22606, new_n22607, new_n22608, new_n22609,
    new_n22611, new_n22612, new_n22613, new_n22614, new_n22615, new_n22616,
    new_n22617, new_n22618, new_n22619, new_n22620, new_n22621, new_n22622,
    new_n22623, new_n22624, new_n22625, new_n22626, new_n22627, new_n22628,
    new_n22629, new_n22630, new_n22631, new_n22632, new_n22633, new_n22634,
    new_n22635, new_n22636, new_n22637, new_n22638, new_n22639, new_n22640,
    new_n22641, new_n22642, new_n22643, new_n22644, new_n22645, new_n22646,
    new_n22647, new_n22648, new_n22649, new_n22650, new_n22651, new_n22652,
    new_n22653, new_n22654, new_n22655, new_n22656, new_n22657, new_n22658,
    new_n22659, new_n22660, new_n22661, new_n22662, new_n22663, new_n22664,
    new_n22665, new_n22666, new_n22667, new_n22668, new_n22669, new_n22670,
    new_n22671, new_n22672, new_n22673, new_n22674, new_n22675, new_n22676,
    new_n22677, new_n22678, new_n22679, new_n22680, new_n22681, new_n22682,
    new_n22683, new_n22684, new_n22685, new_n22686, new_n22687, new_n22688,
    new_n22689, new_n22690, new_n22691, new_n22692, new_n22693, new_n22694,
    new_n22695, new_n22696, new_n22697, new_n22699, new_n22700, new_n22701,
    new_n22702, new_n22703, new_n22704, new_n22705, new_n22706, new_n22707,
    new_n22708, new_n22709, new_n22710, new_n22711, new_n22712, new_n22713,
    new_n22714, new_n22715, new_n22716, new_n22717, new_n22718, new_n22719,
    new_n22720, new_n22721, new_n22722, new_n22723, new_n22724, new_n22725,
    new_n22726, new_n22727, new_n22728, new_n22729, new_n22730, new_n22731,
    new_n22732, new_n22733, new_n22734, new_n22735, new_n22736, new_n22737,
    new_n22738, new_n22739, new_n22740, new_n22741, new_n22742, new_n22743,
    new_n22744, new_n22745, new_n22746, new_n22747, new_n22748, new_n22749,
    new_n22750, new_n22751, new_n22752, new_n22753, new_n22754, new_n22755,
    new_n22756, new_n22757, new_n22758, new_n22759, new_n22760, new_n22761,
    new_n22762, new_n22763, new_n22764, new_n22765, new_n22766, new_n22767,
    new_n22768, new_n22769, new_n22770, new_n22771, new_n22772, new_n22773,
    new_n22774, new_n22775, new_n22776, new_n22777, new_n22778, new_n22779,
    new_n22781, new_n22782, new_n22783, new_n22784, new_n22785, new_n22786,
    new_n22787, new_n22788, new_n22789, new_n22790, new_n22791, new_n22792,
    new_n22793, new_n22794, new_n22795, new_n22796, new_n22797, new_n22798,
    new_n22799, new_n22800, new_n22801, new_n22802, new_n22803, new_n22804,
    new_n22805, new_n22806, new_n22807, new_n22808, new_n22809, new_n22810,
    new_n22811, new_n22812, new_n22813, new_n22814, new_n22815, new_n22816,
    new_n22817, new_n22818, new_n22819, new_n22820, new_n22821, new_n22822,
    new_n22823, new_n22824, new_n22825, new_n22826, new_n22827, new_n22828,
    new_n22829, new_n22830, new_n22831, new_n22832, new_n22833, new_n22834,
    new_n22835, new_n22836, new_n22837, new_n22838, new_n22839, new_n22840,
    new_n22841, new_n22842, new_n22843, new_n22844, new_n22845, new_n22846,
    new_n22847, new_n22848, new_n22849, new_n22850, new_n22851, new_n22852,
    new_n22853, new_n22854, new_n22855, new_n22856, new_n22857, new_n22858,
    new_n22860, new_n22861, new_n22862, new_n22863, new_n22864, new_n22865,
    new_n22866, new_n22867, new_n22868, new_n22869, new_n22870, new_n22871,
    new_n22872, new_n22873, new_n22874, new_n22875, new_n22876, new_n22877,
    new_n22878, new_n22879, new_n22880, new_n22881, new_n22882, new_n22883,
    new_n22884, new_n22885, new_n22886, new_n22887, new_n22888, new_n22889,
    new_n22890, new_n22891, new_n22892, new_n22893, new_n22894, new_n22895,
    new_n22896, new_n22897, new_n22898, new_n22899, new_n22900, new_n22901,
    new_n22902, new_n22903, new_n22904, new_n22905, new_n22906, new_n22907,
    new_n22908, new_n22909, new_n22910, new_n22911, new_n22912, new_n22913,
    new_n22914, new_n22915, new_n22916, new_n22917, new_n22918, new_n22919,
    new_n22920, new_n22921, new_n22922, new_n22923, new_n22924, new_n22925,
    new_n22926, new_n22927, new_n22928, new_n22929, new_n22930, new_n22932,
    new_n22933, new_n22934, new_n22935, new_n22936, new_n22937, new_n22938,
    new_n22939, new_n22940, new_n22941, new_n22942, new_n22943, new_n22944,
    new_n22945, new_n22946, new_n22947, new_n22948, new_n22949, new_n22950,
    new_n22951, new_n22952, new_n22953, new_n22954, new_n22955, new_n22956,
    new_n22957, new_n22958, new_n22959, new_n22960, new_n22961, new_n22962,
    new_n22963, new_n22964, new_n22965, new_n22966, new_n22967, new_n22968,
    new_n22969, new_n22970, new_n22971, new_n22972, new_n22973, new_n22974,
    new_n22975, new_n22976, new_n22977, new_n22978, new_n22979, new_n22980,
    new_n22981, new_n22982, new_n22983, new_n22984, new_n22985, new_n22986,
    new_n22987, new_n22988, new_n22989, new_n22990, new_n22991, new_n22992,
    new_n22993, new_n22994, new_n22995, new_n22997, new_n22998, new_n22999,
    new_n23000, new_n23001, new_n23002, new_n23003, new_n23004, new_n23005,
    new_n23006, new_n23007, new_n23008, new_n23009, new_n23010, new_n23011,
    new_n23012, new_n23013, new_n23014, new_n23015, new_n23016, new_n23017,
    new_n23018, new_n23019, new_n23020, new_n23021, new_n23022, new_n23023,
    new_n23024, new_n23025, new_n23026, new_n23027, new_n23028, new_n23029,
    new_n23030, new_n23031, new_n23032, new_n23033, new_n23034, new_n23035,
    new_n23036, new_n23037, new_n23038, new_n23039, new_n23040, new_n23041,
    new_n23042, new_n23043, new_n23044, new_n23045, new_n23046, new_n23047,
    new_n23048, new_n23049, new_n23050, new_n23051, new_n23052, new_n23053,
    new_n23054, new_n23055, new_n23056, new_n23058, new_n23059, new_n23060,
    new_n23061, new_n23062, new_n23063, new_n23064, new_n23065, new_n23066,
    new_n23067, new_n23068, new_n23069, new_n23070, new_n23071, new_n23072,
    new_n23073, new_n23074, new_n23075, new_n23076, new_n23077, new_n23078,
    new_n23079, new_n23080, new_n23081, new_n23082, new_n23083, new_n23084,
    new_n23085, new_n23086, new_n23087, new_n23088, new_n23089, new_n23090,
    new_n23091, new_n23092, new_n23093, new_n23094, new_n23095, new_n23096,
    new_n23097, new_n23098, new_n23099, new_n23100, new_n23101, new_n23102,
    new_n23103, new_n23104, new_n23105, new_n23106, new_n23107, new_n23108,
    new_n23109, new_n23111, new_n23112, new_n23113, new_n23114, new_n23115,
    new_n23116, new_n23117, new_n23118, new_n23119, new_n23120, new_n23121,
    new_n23122, new_n23123, new_n23124, new_n23125, new_n23126, new_n23127,
    new_n23128, new_n23129, new_n23130, new_n23131, new_n23132, new_n23133,
    new_n23134, new_n23135, new_n23136, new_n23137, new_n23138, new_n23139,
    new_n23140, new_n23141, new_n23142, new_n23143, new_n23144, new_n23145,
    new_n23146, new_n23147, new_n23148, new_n23149, new_n23150, new_n23151,
    new_n23152, new_n23153, new_n23154, new_n23155, new_n23156, new_n23157,
    new_n23158, new_n23160, new_n23161, new_n23162, new_n23163, new_n23164,
    new_n23165, new_n23166, new_n23167, new_n23168, new_n23169, new_n23170,
    new_n23171, new_n23172, new_n23173, new_n23174, new_n23175, new_n23176,
    new_n23177, new_n23178, new_n23179, new_n23180, new_n23181, new_n23182,
    new_n23183, new_n23184, new_n23185, new_n23186, new_n23187, new_n23188,
    new_n23189, new_n23190, new_n23191, new_n23192, new_n23193, new_n23194,
    new_n23195, new_n23196, new_n23197, new_n23198, new_n23199, new_n23200,
    new_n23201, new_n23203, new_n23204, new_n23205, new_n23206, new_n23207,
    new_n23208, new_n23209, new_n23210, new_n23211, new_n23212, new_n23213,
    new_n23214, new_n23215, new_n23216, new_n23217, new_n23218, new_n23219,
    new_n23220, new_n23221, new_n23222, new_n23223, new_n23224, new_n23225,
    new_n23226, new_n23227, new_n23228, new_n23229, new_n23230, new_n23231,
    new_n23232, new_n23233, new_n23234, new_n23235, new_n23236, new_n23237,
    new_n23238, new_n23240, new_n23241, new_n23242, new_n23243, new_n23244,
    new_n23245, new_n23246, new_n23247, new_n23248, new_n23249, new_n23250,
    new_n23251, new_n23252, new_n23253, new_n23254, new_n23255, new_n23256,
    new_n23257, new_n23258, new_n23259, new_n23260, new_n23261, new_n23262,
    new_n23263, new_n23264, new_n23265, new_n23267, new_n23268, new_n23269,
    new_n23270, new_n23271, new_n23272, new_n23273, new_n23274, new_n23275,
    new_n23276, new_n23277, new_n23278, new_n23279, new_n23280, new_n23281,
    new_n23282, new_n23283, new_n23284, new_n23285, new_n23286, new_n23287,
    new_n23288, new_n23289, new_n23290, new_n23292, new_n23293, new_n23294,
    new_n23295, new_n23296, new_n23297, new_n23298, new_n23299, new_n23300,
    new_n23301, new_n23302, new_n23303, new_n23304, new_n23305, new_n23306,
    new_n23307, new_n23309, new_n23310, new_n23311, new_n23312, new_n23313,
    new_n23314, new_n23315, new_n23316, new_n23317, new_n23318, new_n23319,
    new_n23321, new_n23322, new_n23323, new_n23324, new_n23325, new_n23326,
    new_n23327, new_n23329;
  inv1 g00000(.a(\a[1] ), .O(new_n194));
  nor2 g00001(.a(new_n194), .b(\a[0] ), .O(\asquared[2] ));
  inv1 g00002(.a(\a[2] ), .O(new_n196));
  nor2 g00003(.a(new_n196), .b(new_n194), .O(new_n197));
  inv1 g00004(.a(\a[0] ), .O(new_n198));
  nor2 g00005(.a(\a[2] ), .b(\a[1] ), .O(new_n199));
  nor2 g00006(.a(new_n199), .b(new_n198), .O(new_n200));
  inv1 g00007(.a(new_n200), .O(new_n201));
  nor2 g00008(.a(new_n201), .b(new_n197), .O(\asquared[3] ));
  inv1 g00009(.a(\a[3] ), .O(new_n203));
  nor2 g00010(.a(new_n203), .b(new_n196), .O(new_n204));
  inv1 g00011(.a(new_n204), .O(new_n205));
  nor2 g00012(.a(new_n205), .b(new_n198), .O(new_n206));
  nor2 g00013(.a(new_n203), .b(new_n198), .O(new_n207));
  nor2 g00014(.a(\asquared[2] ), .b(new_n196), .O(new_n208));
  nor2 g00015(.a(new_n208), .b(new_n207), .O(new_n209));
  nor2 g00016(.a(new_n209), .b(new_n206), .O(\asquared[4] ));
  inv1 g00017(.a(new_n206), .O(new_n211));
  nor2 g00018(.a(new_n203), .b(new_n194), .O(new_n212));
  inv1 g00019(.a(new_n212), .O(new_n213));
  inv1 g00020(.a(\a[4] ), .O(new_n214));
  nor2 g00021(.a(new_n214), .b(new_n198), .O(new_n215));
  nor2 g00022(.a(new_n215), .b(new_n213), .O(new_n216));
  inv1 g00023(.a(new_n215), .O(new_n217));
  nor2 g00024(.a(new_n217), .b(new_n212), .O(new_n218));
  nor2 g00025(.a(new_n218), .b(new_n216), .O(new_n219));
  inv1 g00026(.a(new_n219), .O(new_n220));
  nor2 g00027(.a(new_n220), .b(new_n197), .O(new_n221));
  inv1 g00028(.a(new_n197), .O(new_n222));
  nor2 g00029(.a(new_n219), .b(new_n222), .O(new_n223));
  nor2 g00030(.a(new_n223), .b(new_n221), .O(new_n224));
  inv1 g00031(.a(new_n224), .O(new_n225));
  nor2 g00032(.a(new_n225), .b(new_n211), .O(new_n226));
  nor2 g00033(.a(new_n224), .b(new_n206), .O(new_n227));
  nor2 g00034(.a(new_n227), .b(new_n226), .O(\asquared[5] ));
  inv1 g00035(.a(\a[5] ), .O(new_n229));
  nor2 g00036(.a(new_n229), .b(new_n198), .O(new_n230));
  inv1 g00037(.a(new_n230), .O(new_n231));
  nor2 g00038(.a(new_n214), .b(new_n194), .O(new_n232));
  inv1 g00039(.a(new_n232), .O(new_n233));
  nor2 g00040(.a(new_n233), .b(new_n207), .O(new_n234));
  nor2 g00041(.a(new_n234), .b(new_n231), .O(new_n235));
  inv1 g00042(.a(new_n234), .O(new_n236));
  nor2 g00043(.a(new_n236), .b(new_n230), .O(new_n237));
  nor2 g00044(.a(new_n237), .b(new_n235), .O(new_n238));
  nor2 g00045(.a(new_n221), .b(new_n211), .O(new_n239));
  nor2 g00046(.a(new_n203), .b(\a[2] ), .O(new_n240));
  nor2 g00047(.a(new_n240), .b(new_n223), .O(new_n241));
  inv1 g00048(.a(new_n241), .O(new_n242));
  nor2 g00049(.a(new_n242), .b(new_n239), .O(new_n243));
  nor2 g00050(.a(new_n243), .b(new_n238), .O(new_n244));
  inv1 g00051(.a(new_n238), .O(new_n245));
  inv1 g00052(.a(new_n243), .O(new_n246));
  nor2 g00053(.a(new_n246), .b(new_n245), .O(new_n247));
  nor2 g00054(.a(new_n247), .b(new_n244), .O(\asquared[6] ));
  inv1 g00055(.a(new_n244), .O(new_n249));
  nor2 g00056(.a(new_n229), .b(new_n194), .O(new_n250));
  nor2 g00057(.a(new_n214), .b(new_n196), .O(new_n251));
  nor2 g00058(.a(new_n251), .b(new_n250), .O(new_n252));
  nor2 g00059(.a(new_n229), .b(new_n196), .O(new_n253));
  inv1 g00060(.a(new_n253), .O(new_n254));
  nor2 g00061(.a(new_n254), .b(new_n233), .O(new_n255));
  nor2 g00062(.a(new_n255), .b(new_n252), .O(new_n256));
  inv1 g00063(.a(\a[6] ), .O(new_n257));
  nor2 g00064(.a(new_n257), .b(new_n198), .O(new_n258));
  nor2 g00065(.a(new_n258), .b(new_n204), .O(new_n259));
  inv1 g00066(.a(new_n207), .O(new_n260));
  nor2 g00067(.a(new_n257), .b(new_n196), .O(new_n261));
  inv1 g00068(.a(new_n261), .O(new_n262));
  nor2 g00069(.a(new_n262), .b(new_n260), .O(new_n263));
  nor2 g00070(.a(new_n263), .b(new_n259), .O(new_n264));
  nor2 g00071(.a(new_n264), .b(new_n256), .O(new_n265));
  inv1 g00072(.a(new_n256), .O(new_n266));
  inv1 g00073(.a(new_n264), .O(new_n267));
  nor2 g00074(.a(new_n267), .b(new_n266), .O(new_n268));
  nor2 g00075(.a(new_n268), .b(new_n265), .O(new_n269));
  nor2 g00076(.a(new_n237), .b(new_n233), .O(new_n270));
  nor2 g00077(.a(new_n270), .b(new_n269), .O(new_n271));
  inv1 g00078(.a(new_n269), .O(new_n272));
  inv1 g00079(.a(new_n270), .O(new_n273));
  nor2 g00080(.a(new_n273), .b(new_n272), .O(new_n274));
  nor2 g00081(.a(new_n274), .b(new_n271), .O(new_n275));
  inv1 g00082(.a(new_n275), .O(new_n276));
  nor2 g00083(.a(new_n276), .b(new_n249), .O(new_n277));
  nor2 g00084(.a(new_n275), .b(new_n244), .O(new_n278));
  nor2 g00085(.a(new_n278), .b(new_n277), .O(\asquared[7] ));
  nor2 g00086(.a(new_n268), .b(new_n263), .O(new_n280));
  nor2 g00087(.a(new_n257), .b(new_n194), .O(new_n281));
  nor2 g00088(.a(new_n281), .b(\a[4] ), .O(new_n282));
  inv1 g00089(.a(new_n281), .O(new_n283));
  nor2 g00090(.a(new_n283), .b(new_n214), .O(new_n284));
  nor2 g00091(.a(new_n284), .b(new_n282), .O(new_n285));
  nor2 g00092(.a(new_n285), .b(new_n255), .O(new_n286));
  inv1 g00093(.a(new_n255), .O(new_n287));
  nor2 g00094(.a(new_n287), .b(\a[6] ), .O(new_n288));
  nor2 g00095(.a(new_n288), .b(new_n286), .O(new_n289));
  inv1 g00096(.a(new_n289), .O(new_n290));
  nor2 g00097(.a(new_n290), .b(new_n280), .O(new_n291));
  inv1 g00098(.a(new_n280), .O(new_n292));
  nor2 g00099(.a(new_n289), .b(new_n292), .O(new_n293));
  nor2 g00100(.a(new_n293), .b(new_n291), .O(new_n294));
  inv1 g00101(.a(\a[7] ), .O(new_n295));
  nor2 g00102(.a(new_n295), .b(new_n198), .O(new_n296));
  inv1 g00103(.a(new_n296), .O(new_n297));
  nor2 g00104(.a(new_n214), .b(new_n203), .O(new_n298));
  nor2 g00105(.a(new_n298), .b(new_n253), .O(new_n299));
  inv1 g00106(.a(new_n251), .O(new_n300));
  nor2 g00107(.a(new_n229), .b(new_n203), .O(new_n301));
  inv1 g00108(.a(new_n301), .O(new_n302));
  nor2 g00109(.a(new_n302), .b(new_n300), .O(new_n303));
  nor2 g00110(.a(new_n303), .b(new_n299), .O(new_n304));
  nor2 g00111(.a(new_n304), .b(new_n297), .O(new_n305));
  inv1 g00112(.a(new_n304), .O(new_n306));
  nor2 g00113(.a(new_n306), .b(new_n296), .O(new_n307));
  nor2 g00114(.a(new_n307), .b(new_n305), .O(new_n308));
  inv1 g00115(.a(new_n308), .O(new_n309));
  nor2 g00116(.a(new_n309), .b(new_n294), .O(new_n310));
  inv1 g00117(.a(new_n294), .O(new_n311));
  nor2 g00118(.a(new_n308), .b(new_n311), .O(new_n312));
  nor2 g00119(.a(new_n312), .b(new_n310), .O(new_n313));
  inv1 g00120(.a(new_n313), .O(new_n314));
  nor2 g00121(.a(new_n277), .b(new_n274), .O(new_n315));
  nor2 g00122(.a(new_n315), .b(new_n314), .O(new_n316));
  inv1 g00123(.a(new_n315), .O(new_n317));
  nor2 g00124(.a(new_n317), .b(new_n313), .O(new_n318));
  nor2 g00125(.a(new_n318), .b(new_n316), .O(\asquared[8] ));
  nor2 g00126(.a(new_n291), .b(new_n288), .O(new_n320));
  inv1 g00127(.a(new_n320), .O(new_n321));
  inv1 g00128(.a(\a[8] ), .O(new_n322));
  nor2 g00129(.a(new_n322), .b(new_n198), .O(new_n323));
  nor2 g00130(.a(new_n323), .b(new_n261), .O(new_n324));
  inv1 g00131(.a(new_n258), .O(new_n325));
  nor2 g00132(.a(new_n322), .b(new_n196), .O(new_n326));
  inv1 g00133(.a(new_n326), .O(new_n327));
  nor2 g00134(.a(new_n327), .b(new_n325), .O(new_n328));
  nor2 g00135(.a(new_n328), .b(new_n324), .O(new_n329));
  inv1 g00136(.a(new_n329), .O(new_n330));
  nor2 g00137(.a(new_n330), .b(new_n284), .O(new_n331));
  inv1 g00138(.a(new_n284), .O(new_n332));
  nor2 g00139(.a(new_n329), .b(new_n332), .O(new_n333));
  nor2 g00140(.a(new_n333), .b(new_n331), .O(new_n334));
  nor2 g00141(.a(new_n295), .b(new_n194), .O(new_n335));
  nor2 g00142(.a(new_n335), .b(new_n301), .O(new_n336));
  inv1 g00143(.a(new_n335), .O(new_n337));
  nor2 g00144(.a(new_n337), .b(new_n302), .O(new_n338));
  nor2 g00145(.a(new_n338), .b(new_n336), .O(new_n339));
  inv1 g00146(.a(new_n339), .O(new_n340));
  nor2 g00147(.a(new_n307), .b(new_n299), .O(new_n341));
  inv1 g00148(.a(new_n341), .O(new_n342));
  nor2 g00149(.a(new_n342), .b(new_n340), .O(new_n343));
  nor2 g00150(.a(new_n341), .b(new_n339), .O(new_n344));
  nor2 g00151(.a(new_n344), .b(new_n343), .O(new_n345));
  inv1 g00152(.a(new_n345), .O(new_n346));
  nor2 g00153(.a(new_n346), .b(new_n334), .O(new_n347));
  inv1 g00154(.a(new_n334), .O(new_n348));
  nor2 g00155(.a(new_n345), .b(new_n348), .O(new_n349));
  nor2 g00156(.a(new_n349), .b(new_n347), .O(new_n350));
  nor2 g00157(.a(new_n350), .b(new_n321), .O(new_n351));
  inv1 g00158(.a(new_n350), .O(new_n352));
  nor2 g00159(.a(new_n352), .b(new_n320), .O(new_n353));
  nor2 g00160(.a(new_n353), .b(new_n351), .O(new_n354));
  inv1 g00161(.a(new_n354), .O(new_n355));
  nor2 g00162(.a(new_n316), .b(new_n312), .O(new_n356));
  nor2 g00163(.a(new_n356), .b(new_n355), .O(new_n357));
  inv1 g00164(.a(new_n356), .O(new_n358));
  nor2 g00165(.a(new_n358), .b(new_n354), .O(new_n359));
  nor2 g00166(.a(new_n359), .b(new_n357), .O(\asquared[9] ));
  nor2 g00167(.a(new_n347), .b(new_n343), .O(new_n361));
  inv1 g00168(.a(new_n338), .O(new_n362));
  inv1 g00169(.a(\a[9] ), .O(new_n363));
  nor2 g00170(.a(new_n363), .b(new_n198), .O(new_n364));
  inv1 g00171(.a(new_n364), .O(new_n365));
  nor2 g00172(.a(new_n365), .b(new_n362), .O(new_n366));
  nor2 g00173(.a(new_n364), .b(new_n338), .O(new_n367));
  nor2 g00174(.a(new_n367), .b(new_n366), .O(new_n368));
  inv1 g00175(.a(new_n368), .O(new_n369));
  nor2 g00176(.a(new_n322), .b(new_n229), .O(new_n370));
  inv1 g00177(.a(new_n370), .O(new_n371));
  nor2 g00178(.a(new_n371), .b(new_n194), .O(new_n372));
  nor2 g00179(.a(new_n372), .b(new_n229), .O(new_n373));
  nor2 g00180(.a(\a[5] ), .b(new_n194), .O(new_n374));
  inv1 g00181(.a(new_n374), .O(new_n375));
  nor2 g00182(.a(new_n375), .b(new_n322), .O(new_n376));
  nor2 g00183(.a(new_n376), .b(new_n373), .O(new_n377));
  nor2 g00184(.a(new_n377), .b(new_n369), .O(new_n378));
  inv1 g00185(.a(new_n377), .O(new_n379));
  nor2 g00186(.a(new_n379), .b(new_n368), .O(new_n380));
  nor2 g00187(.a(new_n380), .b(new_n378), .O(new_n381));
  inv1 g00188(.a(new_n381), .O(new_n382));
  nor2 g00189(.a(new_n295), .b(new_n196), .O(new_n383));
  nor2 g00190(.a(new_n229), .b(new_n214), .O(new_n384));
  nor2 g00191(.a(new_n257), .b(new_n203), .O(new_n385));
  nor2 g00192(.a(new_n385), .b(new_n384), .O(new_n386));
  nor2 g00193(.a(new_n257), .b(new_n214), .O(new_n387));
  inv1 g00194(.a(new_n387), .O(new_n388));
  nor2 g00195(.a(new_n388), .b(new_n302), .O(new_n389));
  nor2 g00196(.a(new_n389), .b(new_n386), .O(new_n390));
  inv1 g00197(.a(new_n390), .O(new_n391));
  nor2 g00198(.a(new_n391), .b(new_n383), .O(new_n392));
  inv1 g00199(.a(new_n383), .O(new_n393));
  nor2 g00200(.a(new_n390), .b(new_n393), .O(new_n394));
  nor2 g00201(.a(new_n394), .b(new_n392), .O(new_n395));
  nor2 g00202(.a(new_n331), .b(new_n324), .O(new_n396));
  inv1 g00203(.a(new_n396), .O(new_n397));
  nor2 g00204(.a(new_n397), .b(new_n395), .O(new_n398));
  inv1 g00205(.a(new_n395), .O(new_n399));
  nor2 g00206(.a(new_n396), .b(new_n399), .O(new_n400));
  nor2 g00207(.a(new_n400), .b(new_n398), .O(new_n401));
  inv1 g00208(.a(new_n401), .O(new_n402));
  nor2 g00209(.a(new_n402), .b(new_n382), .O(new_n403));
  nor2 g00210(.a(new_n401), .b(new_n381), .O(new_n404));
  nor2 g00211(.a(new_n404), .b(new_n403), .O(new_n405));
  inv1 g00212(.a(new_n405), .O(new_n406));
  nor2 g00213(.a(new_n406), .b(new_n361), .O(new_n407));
  inv1 g00214(.a(new_n361), .O(new_n408));
  nor2 g00215(.a(new_n405), .b(new_n408), .O(new_n409));
  nor2 g00216(.a(new_n409), .b(new_n407), .O(new_n410));
  inv1 g00217(.a(new_n410), .O(new_n411));
  nor2 g00218(.a(new_n357), .b(new_n353), .O(new_n412));
  nor2 g00219(.a(new_n412), .b(new_n411), .O(new_n413));
  inv1 g00220(.a(new_n412), .O(new_n414));
  nor2 g00221(.a(new_n414), .b(new_n410), .O(new_n415));
  nor2 g00222(.a(new_n415), .b(new_n413), .O(\asquared[10] ));
  nor2 g00223(.a(new_n403), .b(new_n398), .O(new_n417));
  inv1 g00224(.a(new_n417), .O(new_n418));
  inv1 g00225(.a(new_n372), .O(new_n419));
  nor2 g00226(.a(new_n363), .b(new_n194), .O(new_n420));
  nor2 g00227(.a(new_n420), .b(new_n387), .O(new_n421));
  nor2 g00228(.a(new_n363), .b(new_n214), .O(new_n422));
  inv1 g00229(.a(new_n422), .O(new_n423));
  nor2 g00230(.a(new_n423), .b(new_n283), .O(new_n424));
  nor2 g00231(.a(new_n424), .b(new_n421), .O(new_n425));
  inv1 g00232(.a(new_n425), .O(new_n426));
  nor2 g00233(.a(new_n426), .b(new_n419), .O(new_n427));
  nor2 g00234(.a(new_n425), .b(new_n372), .O(new_n428));
  nor2 g00235(.a(new_n428), .b(new_n427), .O(new_n429));
  inv1 g00236(.a(new_n429), .O(new_n430));
  nor2 g00237(.a(new_n392), .b(new_n386), .O(new_n431));
  inv1 g00238(.a(new_n431), .O(new_n432));
  nor2 g00239(.a(new_n432), .b(new_n430), .O(new_n433));
  nor2 g00240(.a(new_n431), .b(new_n429), .O(new_n434));
  nor2 g00241(.a(new_n434), .b(new_n433), .O(new_n435));
  inv1 g00242(.a(new_n435), .O(new_n436));
  nor2 g00243(.a(new_n295), .b(new_n203), .O(new_n437));
  inv1 g00244(.a(\a[10] ), .O(new_n438));
  nor2 g00245(.a(new_n438), .b(new_n198), .O(new_n439));
  nor2 g00246(.a(new_n439), .b(new_n437), .O(new_n440));
  inv1 g00247(.a(new_n437), .O(new_n441));
  inv1 g00248(.a(new_n439), .O(new_n442));
  nor2 g00249(.a(new_n442), .b(new_n441), .O(new_n443));
  nor2 g00250(.a(new_n443), .b(new_n440), .O(new_n444));
  nor2 g00251(.a(new_n444), .b(new_n327), .O(new_n445));
  inv1 g00252(.a(new_n444), .O(new_n446));
  nor2 g00253(.a(new_n446), .b(new_n326), .O(new_n447));
  nor2 g00254(.a(new_n447), .b(new_n445), .O(new_n448));
  nor2 g00255(.a(new_n378), .b(new_n366), .O(new_n449));
  nor2 g00256(.a(new_n449), .b(new_n448), .O(new_n450));
  inv1 g00257(.a(new_n448), .O(new_n451));
  inv1 g00258(.a(new_n449), .O(new_n452));
  nor2 g00259(.a(new_n452), .b(new_n451), .O(new_n453));
  nor2 g00260(.a(new_n453), .b(new_n450), .O(new_n454));
  inv1 g00261(.a(new_n454), .O(new_n455));
  nor2 g00262(.a(new_n455), .b(new_n436), .O(new_n456));
  nor2 g00263(.a(new_n454), .b(new_n435), .O(new_n457));
  nor2 g00264(.a(new_n457), .b(new_n456), .O(new_n458));
  nor2 g00265(.a(new_n458), .b(new_n418), .O(new_n459));
  inv1 g00266(.a(new_n458), .O(new_n460));
  nor2 g00267(.a(new_n460), .b(new_n417), .O(new_n461));
  nor2 g00268(.a(new_n461), .b(new_n459), .O(new_n462));
  inv1 g00269(.a(new_n462), .O(new_n463));
  nor2 g00270(.a(new_n413), .b(new_n407), .O(new_n464));
  nor2 g00271(.a(new_n464), .b(new_n463), .O(new_n465));
  inv1 g00272(.a(new_n464), .O(new_n466));
  nor2 g00273(.a(new_n466), .b(new_n462), .O(new_n467));
  nor2 g00274(.a(new_n467), .b(new_n465), .O(\asquared[11] ));
  nor2 g00275(.a(new_n456), .b(new_n450), .O(new_n469));
  inv1 g00276(.a(new_n469), .O(new_n470));
  inv1 g00277(.a(new_n424), .O(new_n471));
  nor2 g00278(.a(new_n363), .b(new_n196), .O(new_n472));
  nor2 g00279(.a(new_n322), .b(new_n203), .O(new_n473));
  nor2 g00280(.a(new_n473), .b(new_n472), .O(new_n474));
  nor2 g00281(.a(new_n363), .b(new_n203), .O(new_n475));
  inv1 g00282(.a(new_n475), .O(new_n476));
  nor2 g00283(.a(new_n476), .b(new_n327), .O(new_n477));
  nor2 g00284(.a(new_n477), .b(new_n474), .O(new_n478));
  nor2 g00285(.a(new_n478), .b(new_n471), .O(new_n479));
  inv1 g00286(.a(new_n478), .O(new_n480));
  nor2 g00287(.a(new_n480), .b(new_n424), .O(new_n481));
  nor2 g00288(.a(new_n481), .b(new_n479), .O(new_n482));
  nor2 g00289(.a(new_n283), .b(new_n438), .O(new_n483));
  nor2 g00290(.a(new_n483), .b(new_n257), .O(new_n484));
  nor2 g00291(.a(\a[6] ), .b(new_n194), .O(new_n485));
  inv1 g00292(.a(new_n485), .O(new_n486));
  nor2 g00293(.a(new_n486), .b(new_n438), .O(new_n487));
  nor2 g00294(.a(new_n487), .b(new_n484), .O(new_n488));
  nor2 g00295(.a(new_n447), .b(new_n440), .O(new_n489));
  inv1 g00296(.a(new_n489), .O(new_n490));
  nor2 g00297(.a(new_n490), .b(new_n488), .O(new_n491));
  inv1 g00298(.a(new_n488), .O(new_n492));
  nor2 g00299(.a(new_n489), .b(new_n492), .O(new_n493));
  nor2 g00300(.a(new_n493), .b(new_n491), .O(new_n494));
  inv1 g00301(.a(new_n494), .O(new_n495));
  nor2 g00302(.a(new_n495), .b(new_n482), .O(new_n496));
  inv1 g00303(.a(new_n482), .O(new_n497));
  nor2 g00304(.a(new_n494), .b(new_n497), .O(new_n498));
  nor2 g00305(.a(new_n498), .b(new_n496), .O(new_n499));
  inv1 g00306(.a(new_n499), .O(new_n500));
  nor2 g00307(.a(new_n433), .b(new_n427), .O(new_n501));
  inv1 g00308(.a(\a[11] ), .O(new_n502));
  nor2 g00309(.a(new_n502), .b(new_n198), .O(new_n503));
  nor2 g00310(.a(new_n257), .b(new_n229), .O(new_n504));
  nor2 g00311(.a(new_n295), .b(new_n214), .O(new_n505));
  nor2 g00312(.a(new_n505), .b(new_n504), .O(new_n506));
  nor2 g00313(.a(new_n295), .b(new_n229), .O(new_n507));
  inv1 g00314(.a(new_n507), .O(new_n508));
  nor2 g00315(.a(new_n508), .b(new_n388), .O(new_n509));
  nor2 g00316(.a(new_n509), .b(new_n506), .O(new_n510));
  inv1 g00317(.a(new_n510), .O(new_n511));
  nor2 g00318(.a(new_n511), .b(new_n503), .O(new_n512));
  inv1 g00319(.a(new_n503), .O(new_n513));
  nor2 g00320(.a(new_n510), .b(new_n513), .O(new_n514));
  nor2 g00321(.a(new_n514), .b(new_n512), .O(new_n515));
  nor2 g00322(.a(new_n515), .b(new_n501), .O(new_n516));
  inv1 g00323(.a(new_n501), .O(new_n517));
  inv1 g00324(.a(new_n515), .O(new_n518));
  nor2 g00325(.a(new_n518), .b(new_n517), .O(new_n519));
  nor2 g00326(.a(new_n519), .b(new_n516), .O(new_n520));
  inv1 g00327(.a(new_n520), .O(new_n521));
  nor2 g00328(.a(new_n521), .b(new_n500), .O(new_n522));
  nor2 g00329(.a(new_n520), .b(new_n499), .O(new_n523));
  nor2 g00330(.a(new_n523), .b(new_n522), .O(new_n524));
  nor2 g00331(.a(new_n524), .b(new_n470), .O(new_n525));
  inv1 g00332(.a(new_n524), .O(new_n526));
  nor2 g00333(.a(new_n526), .b(new_n469), .O(new_n527));
  nor2 g00334(.a(new_n527), .b(new_n525), .O(new_n528));
  inv1 g00335(.a(new_n528), .O(new_n529));
  nor2 g00336(.a(new_n465), .b(new_n461), .O(new_n530));
  nor2 g00337(.a(new_n530), .b(new_n529), .O(new_n531));
  inv1 g00338(.a(new_n530), .O(new_n532));
  nor2 g00339(.a(new_n532), .b(new_n528), .O(new_n533));
  nor2 g00340(.a(new_n533), .b(new_n531), .O(\asquared[12] ));
  nor2 g00341(.a(new_n522), .b(new_n516), .O(new_n535));
  inv1 g00342(.a(new_n535), .O(new_n536));
  nor2 g00343(.a(new_n496), .b(new_n491), .O(new_n537));
  nor2 g00344(.a(new_n502), .b(new_n194), .O(new_n538));
  nor2 g00345(.a(new_n538), .b(new_n507), .O(new_n539));
  nor2 g00346(.a(new_n502), .b(new_n229), .O(new_n540));
  inv1 g00347(.a(new_n540), .O(new_n541));
  nor2 g00348(.a(new_n541), .b(new_n337), .O(new_n542));
  nor2 g00349(.a(new_n542), .b(new_n539), .O(new_n543));
  inv1 g00350(.a(new_n543), .O(new_n544));
  nor2 g00351(.a(new_n322), .b(new_n214), .O(new_n545));
  nor2 g00352(.a(new_n545), .b(new_n483), .O(new_n546));
  inv1 g00353(.a(new_n483), .O(new_n547));
  inv1 g00354(.a(new_n545), .O(new_n548));
  nor2 g00355(.a(new_n548), .b(new_n547), .O(new_n549));
  nor2 g00356(.a(new_n549), .b(new_n546), .O(new_n550));
  nor2 g00357(.a(new_n550), .b(new_n544), .O(new_n551));
  inv1 g00358(.a(new_n550), .O(new_n552));
  nor2 g00359(.a(new_n552), .b(new_n543), .O(new_n553));
  nor2 g00360(.a(new_n553), .b(new_n551), .O(new_n554));
  nor2 g00361(.a(new_n554), .b(new_n537), .O(new_n555));
  inv1 g00362(.a(new_n537), .O(new_n556));
  inv1 g00363(.a(new_n554), .O(new_n557));
  nor2 g00364(.a(new_n557), .b(new_n556), .O(new_n558));
  nor2 g00365(.a(new_n558), .b(new_n555), .O(new_n559));
  inv1 g00366(.a(new_n559), .O(new_n560));
  nor2 g00367(.a(new_n481), .b(new_n474), .O(new_n561));
  nor2 g00368(.a(new_n512), .b(new_n506), .O(new_n562));
  nor2 g00369(.a(new_n562), .b(new_n561), .O(new_n563));
  inv1 g00370(.a(new_n561), .O(new_n564));
  inv1 g00371(.a(new_n562), .O(new_n565));
  nor2 g00372(.a(new_n565), .b(new_n564), .O(new_n566));
  nor2 g00373(.a(new_n566), .b(new_n563), .O(new_n567));
  inv1 g00374(.a(new_n567), .O(new_n568));
  inv1 g00375(.a(\a[12] ), .O(new_n569));
  nor2 g00376(.a(new_n569), .b(new_n198), .O(new_n570));
  nor2 g00377(.a(new_n438), .b(new_n196), .O(new_n571));
  nor2 g00378(.a(new_n571), .b(new_n570), .O(new_n572));
  nor2 g00379(.a(new_n569), .b(new_n196), .O(new_n573));
  inv1 g00380(.a(new_n573), .O(new_n574));
  nor2 g00381(.a(new_n574), .b(new_n442), .O(new_n575));
  nor2 g00382(.a(new_n575), .b(new_n572), .O(new_n576));
  nor2 g00383(.a(new_n576), .b(new_n476), .O(new_n577));
  inv1 g00384(.a(new_n576), .O(new_n578));
  nor2 g00385(.a(new_n578), .b(new_n475), .O(new_n579));
  nor2 g00386(.a(new_n579), .b(new_n577), .O(new_n580));
  inv1 g00387(.a(new_n580), .O(new_n581));
  nor2 g00388(.a(new_n581), .b(new_n568), .O(new_n582));
  nor2 g00389(.a(new_n580), .b(new_n567), .O(new_n583));
  nor2 g00390(.a(new_n583), .b(new_n582), .O(new_n584));
  nor2 g00391(.a(new_n584), .b(new_n560), .O(new_n585));
  inv1 g00392(.a(new_n584), .O(new_n586));
  nor2 g00393(.a(new_n586), .b(new_n559), .O(new_n587));
  nor2 g00394(.a(new_n587), .b(new_n585), .O(new_n588));
  nor2 g00395(.a(new_n588), .b(new_n536), .O(new_n589));
  inv1 g00396(.a(new_n588), .O(new_n590));
  nor2 g00397(.a(new_n590), .b(new_n535), .O(new_n591));
  nor2 g00398(.a(new_n591), .b(new_n589), .O(new_n592));
  inv1 g00399(.a(new_n592), .O(new_n593));
  nor2 g00400(.a(new_n531), .b(new_n527), .O(new_n594));
  nor2 g00401(.a(new_n594), .b(new_n593), .O(new_n595));
  inv1 g00402(.a(new_n594), .O(new_n596));
  nor2 g00403(.a(new_n596), .b(new_n592), .O(new_n597));
  nor2 g00404(.a(new_n597), .b(new_n595), .O(\asquared[13] ));
  nor2 g00405(.a(new_n502), .b(new_n196), .O(new_n599));
  inv1 g00406(.a(new_n599), .O(new_n600));
  nor2 g00407(.a(new_n295), .b(new_n257), .O(new_n601));
  nor2 g00408(.a(new_n601), .b(new_n370), .O(new_n602));
  nor2 g00409(.a(new_n322), .b(new_n257), .O(new_n603));
  inv1 g00410(.a(new_n603), .O(new_n604));
  nor2 g00411(.a(new_n604), .b(new_n508), .O(new_n605));
  nor2 g00412(.a(new_n605), .b(new_n602), .O(new_n606));
  nor2 g00413(.a(new_n606), .b(new_n600), .O(new_n607));
  inv1 g00414(.a(new_n606), .O(new_n608));
  nor2 g00415(.a(new_n608), .b(new_n599), .O(new_n609));
  nor2 g00416(.a(new_n609), .b(new_n607), .O(new_n610));
  nor2 g00417(.a(new_n438), .b(new_n203), .O(new_n611));
  inv1 g00418(.a(new_n611), .O(new_n612));
  inv1 g00419(.a(\a[13] ), .O(new_n613));
  nor2 g00420(.a(new_n613), .b(new_n198), .O(new_n614));
  nor2 g00421(.a(new_n614), .b(new_n422), .O(new_n615));
  nor2 g00422(.a(new_n613), .b(new_n214), .O(new_n616));
  inv1 g00423(.a(new_n616), .O(new_n617));
  nor2 g00424(.a(new_n617), .b(new_n365), .O(new_n618));
  nor2 g00425(.a(new_n618), .b(new_n615), .O(new_n619));
  nor2 g00426(.a(new_n619), .b(new_n612), .O(new_n620));
  inv1 g00427(.a(new_n619), .O(new_n621));
  nor2 g00428(.a(new_n621), .b(new_n611), .O(new_n622));
  nor2 g00429(.a(new_n622), .b(new_n620), .O(new_n623));
  nor2 g00430(.a(new_n553), .b(new_n546), .O(new_n624));
  inv1 g00431(.a(new_n624), .O(new_n625));
  nor2 g00432(.a(new_n625), .b(new_n623), .O(new_n626));
  inv1 g00433(.a(new_n623), .O(new_n627));
  nor2 g00434(.a(new_n624), .b(new_n627), .O(new_n628));
  nor2 g00435(.a(new_n628), .b(new_n626), .O(new_n629));
  inv1 g00436(.a(new_n629), .O(new_n630));
  nor2 g00437(.a(new_n630), .b(new_n610), .O(new_n631));
  inv1 g00438(.a(new_n610), .O(new_n632));
  nor2 g00439(.a(new_n629), .b(new_n632), .O(new_n633));
  nor2 g00440(.a(new_n633), .b(new_n631), .O(new_n634));
  inv1 g00441(.a(new_n542), .O(new_n635));
  nor2 g00442(.a(new_n635), .b(\a[12] ), .O(new_n636));
  nor2 g00443(.a(new_n337), .b(new_n569), .O(new_n637));
  nor2 g00444(.a(new_n569), .b(new_n194), .O(new_n638));
  nor2 g00445(.a(new_n638), .b(\a[7] ), .O(new_n639));
  nor2 g00446(.a(new_n639), .b(new_n637), .O(new_n640));
  nor2 g00447(.a(new_n640), .b(new_n542), .O(new_n641));
  nor2 g00448(.a(new_n641), .b(new_n636), .O(new_n642));
  inv1 g00449(.a(new_n642), .O(new_n643));
  nor2 g00450(.a(new_n579), .b(new_n572), .O(new_n644));
  inv1 g00451(.a(new_n644), .O(new_n645));
  nor2 g00452(.a(new_n645), .b(new_n643), .O(new_n646));
  nor2 g00453(.a(new_n644), .b(new_n642), .O(new_n647));
  nor2 g00454(.a(new_n647), .b(new_n646), .O(new_n648));
  nor2 g00455(.a(new_n582), .b(new_n563), .O(new_n649));
  nor2 g00456(.a(new_n649), .b(new_n648), .O(new_n650));
  inv1 g00457(.a(new_n648), .O(new_n651));
  inv1 g00458(.a(new_n649), .O(new_n652));
  nor2 g00459(.a(new_n652), .b(new_n651), .O(new_n653));
  nor2 g00460(.a(new_n653), .b(new_n650), .O(new_n654));
  nor2 g00461(.a(new_n585), .b(new_n555), .O(new_n655));
  inv1 g00462(.a(new_n655), .O(new_n656));
  nor2 g00463(.a(new_n656), .b(new_n654), .O(new_n657));
  inv1 g00464(.a(new_n654), .O(new_n658));
  nor2 g00465(.a(new_n655), .b(new_n658), .O(new_n659));
  nor2 g00466(.a(new_n659), .b(new_n657), .O(new_n660));
  nor2 g00467(.a(new_n660), .b(new_n634), .O(new_n661));
  inv1 g00468(.a(new_n634), .O(new_n662));
  inv1 g00469(.a(new_n660), .O(new_n663));
  nor2 g00470(.a(new_n663), .b(new_n662), .O(new_n664));
  nor2 g00471(.a(new_n664), .b(new_n661), .O(new_n665));
  inv1 g00472(.a(new_n665), .O(new_n666));
  nor2 g00473(.a(new_n595), .b(new_n591), .O(new_n667));
  nor2 g00474(.a(new_n667), .b(new_n666), .O(new_n668));
  inv1 g00475(.a(new_n667), .O(new_n669));
  nor2 g00476(.a(new_n669), .b(new_n665), .O(new_n670));
  nor2 g00477(.a(new_n670), .b(new_n668), .O(\asquared[14] ));
  nor2 g00478(.a(new_n659), .b(new_n653), .O(new_n672));
  nor2 g00479(.a(new_n631), .b(new_n626), .O(new_n673));
  inv1 g00480(.a(new_n673), .O(new_n674));
  nor2 g00481(.a(new_n613), .b(new_n194), .O(new_n675));
  nor2 g00482(.a(new_n675), .b(new_n603), .O(new_n676));
  inv1 g00483(.a(new_n675), .O(new_n677));
  nor2 g00484(.a(new_n677), .b(new_n604), .O(new_n678));
  nor2 g00485(.a(new_n678), .b(new_n676), .O(new_n679));
  inv1 g00486(.a(new_n679), .O(new_n680));
  nor2 g00487(.a(new_n609), .b(new_n602), .O(new_n681));
  inv1 g00488(.a(new_n681), .O(new_n682));
  nor2 g00489(.a(new_n682), .b(new_n680), .O(new_n683));
  nor2 g00490(.a(new_n681), .b(new_n679), .O(new_n684));
  nor2 g00491(.a(new_n684), .b(new_n683), .O(new_n685));
  inv1 g00492(.a(new_n685), .O(new_n686));
  nor2 g00493(.a(new_n622), .b(new_n615), .O(new_n687));
  inv1 g00494(.a(new_n687), .O(new_n688));
  nor2 g00495(.a(new_n688), .b(new_n686), .O(new_n689));
  nor2 g00496(.a(new_n687), .b(new_n685), .O(new_n690));
  nor2 g00497(.a(new_n690), .b(new_n689), .O(new_n691));
  nor2 g00498(.a(new_n691), .b(new_n674), .O(new_n692));
  inv1 g00499(.a(new_n691), .O(new_n693));
  nor2 g00500(.a(new_n693), .b(new_n673), .O(new_n694));
  nor2 g00501(.a(new_n694), .b(new_n692), .O(new_n695));
  inv1 g00502(.a(new_n695), .O(new_n696));
  nor2 g00503(.a(new_n646), .b(new_n636), .O(new_n697));
  inv1 g00504(.a(new_n697), .O(new_n698));
  inv1 g00505(.a(\a[14] ), .O(new_n699));
  nor2 g00506(.a(new_n699), .b(new_n198), .O(new_n700));
  nor2 g00507(.a(new_n502), .b(new_n203), .O(new_n701));
  nor2 g00508(.a(new_n701), .b(new_n573), .O(new_n702));
  nor2 g00509(.a(new_n569), .b(new_n203), .O(new_n703));
  inv1 g00510(.a(new_n703), .O(new_n704));
  nor2 g00511(.a(new_n704), .b(new_n600), .O(new_n705));
  nor2 g00512(.a(new_n705), .b(new_n702), .O(new_n706));
  inv1 g00513(.a(new_n706), .O(new_n707));
  nor2 g00514(.a(new_n707), .b(new_n700), .O(new_n708));
  inv1 g00515(.a(new_n700), .O(new_n709));
  nor2 g00516(.a(new_n706), .b(new_n709), .O(new_n710));
  nor2 g00517(.a(new_n710), .b(new_n708), .O(new_n711));
  inv1 g00518(.a(new_n637), .O(new_n712));
  nor2 g00519(.a(new_n438), .b(new_n214), .O(new_n713));
  nor2 g00520(.a(new_n363), .b(new_n229), .O(new_n714));
  nor2 g00521(.a(new_n714), .b(new_n713), .O(new_n715));
  nor2 g00522(.a(new_n438), .b(new_n229), .O(new_n716));
  inv1 g00523(.a(new_n716), .O(new_n717));
  nor2 g00524(.a(new_n717), .b(new_n423), .O(new_n718));
  nor2 g00525(.a(new_n718), .b(new_n715), .O(new_n719));
  nor2 g00526(.a(new_n719), .b(new_n712), .O(new_n720));
  inv1 g00527(.a(new_n719), .O(new_n721));
  nor2 g00528(.a(new_n721), .b(new_n637), .O(new_n722));
  nor2 g00529(.a(new_n722), .b(new_n720), .O(new_n723));
  nor2 g00530(.a(new_n723), .b(new_n711), .O(new_n724));
  inv1 g00531(.a(new_n711), .O(new_n725));
  inv1 g00532(.a(new_n723), .O(new_n726));
  nor2 g00533(.a(new_n726), .b(new_n725), .O(new_n727));
  nor2 g00534(.a(new_n727), .b(new_n724), .O(new_n728));
  nor2 g00535(.a(new_n728), .b(new_n698), .O(new_n729));
  inv1 g00536(.a(new_n728), .O(new_n730));
  nor2 g00537(.a(new_n730), .b(new_n697), .O(new_n731));
  nor2 g00538(.a(new_n731), .b(new_n729), .O(new_n732));
  inv1 g00539(.a(new_n732), .O(new_n733));
  nor2 g00540(.a(new_n733), .b(new_n696), .O(new_n734));
  nor2 g00541(.a(new_n732), .b(new_n695), .O(new_n735));
  nor2 g00542(.a(new_n735), .b(new_n734), .O(new_n736));
  inv1 g00543(.a(new_n736), .O(new_n737));
  nor2 g00544(.a(new_n737), .b(new_n672), .O(new_n738));
  inv1 g00545(.a(new_n672), .O(new_n739));
  nor2 g00546(.a(new_n736), .b(new_n739), .O(new_n740));
  nor2 g00547(.a(new_n740), .b(new_n738), .O(new_n741));
  nor2 g00548(.a(new_n668), .b(new_n664), .O(new_n742));
  inv1 g00549(.a(new_n742), .O(new_n743));
  nor2 g00550(.a(new_n743), .b(new_n741), .O(new_n744));
  inv1 g00551(.a(new_n741), .O(new_n745));
  nor2 g00552(.a(new_n742), .b(new_n745), .O(new_n746));
  nor2 g00553(.a(new_n746), .b(new_n744), .O(\asquared[15] ));
  nor2 g00554(.a(new_n734), .b(new_n694), .O(new_n748));
  nor2 g00555(.a(new_n689), .b(new_n683), .O(new_n749));
  inv1 g00556(.a(new_n749), .O(new_n750));
  nor2 g00557(.a(new_n613), .b(new_n196), .O(new_n751));
  inv1 g00558(.a(new_n751), .O(new_n752));
  nor2 g00559(.a(new_n322), .b(new_n295), .O(new_n753));
  nor2 g00560(.a(new_n363), .b(new_n257), .O(new_n754));
  nor2 g00561(.a(new_n754), .b(new_n753), .O(new_n755));
  inv1 g00562(.a(new_n753), .O(new_n756));
  inv1 g00563(.a(new_n754), .O(new_n757));
  nor2 g00564(.a(new_n757), .b(new_n756), .O(new_n758));
  nor2 g00565(.a(new_n758), .b(new_n755), .O(new_n759));
  nor2 g00566(.a(new_n759), .b(new_n752), .O(new_n760));
  inv1 g00567(.a(new_n759), .O(new_n761));
  nor2 g00568(.a(new_n761), .b(new_n751), .O(new_n762));
  nor2 g00569(.a(new_n762), .b(new_n760), .O(new_n763));
  nor2 g00570(.a(new_n502), .b(new_n214), .O(new_n764));
  nor2 g00571(.a(new_n764), .b(new_n678), .O(new_n765));
  inv1 g00572(.a(new_n678), .O(new_n766));
  inv1 g00573(.a(new_n764), .O(new_n767));
  nor2 g00574(.a(new_n767), .b(new_n766), .O(new_n768));
  nor2 g00575(.a(new_n768), .b(new_n765), .O(new_n769));
  inv1 g00576(.a(new_n769), .O(new_n770));
  nor2 g00577(.a(new_n699), .b(new_n194), .O(new_n771));
  inv1 g00578(.a(new_n771), .O(new_n772));
  nor2 g00579(.a(new_n772), .b(new_n322), .O(new_n773));
  nor2 g00580(.a(new_n771), .b(\a[8] ), .O(new_n774));
  nor2 g00581(.a(new_n774), .b(new_n773), .O(new_n775));
  inv1 g00582(.a(new_n775), .O(new_n776));
  nor2 g00583(.a(new_n776), .b(new_n770), .O(new_n777));
  nor2 g00584(.a(new_n775), .b(new_n769), .O(new_n778));
  nor2 g00585(.a(new_n778), .b(new_n777), .O(new_n779));
  inv1 g00586(.a(new_n779), .O(new_n780));
  nor2 g00587(.a(new_n780), .b(new_n763), .O(new_n781));
  inv1 g00588(.a(new_n763), .O(new_n782));
  nor2 g00589(.a(new_n779), .b(new_n782), .O(new_n783));
  nor2 g00590(.a(new_n783), .b(new_n781), .O(new_n784));
  nor2 g00591(.a(new_n784), .b(new_n750), .O(new_n785));
  inv1 g00592(.a(new_n784), .O(new_n786));
  nor2 g00593(.a(new_n786), .b(new_n749), .O(new_n787));
  nor2 g00594(.a(new_n787), .b(new_n785), .O(new_n788));
  inv1 g00595(.a(new_n788), .O(new_n789));
  nor2 g00596(.a(new_n731), .b(new_n724), .O(new_n790));
  inv1 g00597(.a(new_n790), .O(new_n791));
  nor2 g00598(.a(new_n722), .b(new_n715), .O(new_n792));
  nor2 g00599(.a(new_n708), .b(new_n702), .O(new_n793));
  nor2 g00600(.a(new_n793), .b(new_n792), .O(new_n794));
  inv1 g00601(.a(new_n792), .O(new_n795));
  inv1 g00602(.a(new_n793), .O(new_n796));
  nor2 g00603(.a(new_n796), .b(new_n795), .O(new_n797));
  nor2 g00604(.a(new_n797), .b(new_n794), .O(new_n798));
  inv1 g00605(.a(new_n798), .O(new_n799));
  inv1 g00606(.a(\a[15] ), .O(new_n800));
  nor2 g00607(.a(new_n800), .b(new_n198), .O(new_n801));
  nor2 g00608(.a(new_n801), .b(new_n703), .O(new_n802));
  inv1 g00609(.a(new_n801), .O(new_n803));
  nor2 g00610(.a(new_n803), .b(new_n704), .O(new_n804));
  nor2 g00611(.a(new_n804), .b(new_n802), .O(new_n805));
  nor2 g00612(.a(new_n805), .b(new_n717), .O(new_n806));
  inv1 g00613(.a(new_n805), .O(new_n807));
  nor2 g00614(.a(new_n807), .b(new_n716), .O(new_n808));
  nor2 g00615(.a(new_n808), .b(new_n806), .O(new_n809));
  inv1 g00616(.a(new_n809), .O(new_n810));
  nor2 g00617(.a(new_n810), .b(new_n799), .O(new_n811));
  nor2 g00618(.a(new_n809), .b(new_n798), .O(new_n812));
  nor2 g00619(.a(new_n812), .b(new_n811), .O(new_n813));
  inv1 g00620(.a(new_n813), .O(new_n814));
  nor2 g00621(.a(new_n814), .b(new_n791), .O(new_n815));
  nor2 g00622(.a(new_n813), .b(new_n790), .O(new_n816));
  nor2 g00623(.a(new_n816), .b(new_n815), .O(new_n817));
  inv1 g00624(.a(new_n817), .O(new_n818));
  nor2 g00625(.a(new_n818), .b(new_n789), .O(new_n819));
  nor2 g00626(.a(new_n817), .b(new_n788), .O(new_n820));
  nor2 g00627(.a(new_n820), .b(new_n819), .O(new_n821));
  inv1 g00628(.a(new_n821), .O(new_n822));
  nor2 g00629(.a(new_n822), .b(new_n748), .O(new_n823));
  inv1 g00630(.a(new_n748), .O(new_n824));
  nor2 g00631(.a(new_n821), .b(new_n824), .O(new_n825));
  nor2 g00632(.a(new_n825), .b(new_n823), .O(new_n826));
  inv1 g00633(.a(new_n826), .O(new_n827));
  nor2 g00634(.a(new_n743), .b(new_n738), .O(new_n828));
  nor2 g00635(.a(new_n828), .b(new_n740), .O(new_n829));
  nor2 g00636(.a(new_n829), .b(new_n827), .O(new_n830));
  inv1 g00637(.a(new_n829), .O(new_n831));
  nor2 g00638(.a(new_n831), .b(new_n826), .O(new_n832));
  nor2 g00639(.a(new_n832), .b(new_n830), .O(new_n833));
  inv1 g00640(.a(new_n833), .O(\asquared[16] ));
  nor2 g00641(.a(new_n819), .b(new_n816), .O(new_n835));
  nor2 g00642(.a(new_n787), .b(new_n781), .O(new_n836));
  inv1 g00643(.a(new_n836), .O(new_n837));
  nor2 g00644(.a(new_n777), .b(new_n768), .O(new_n838));
  inv1 g00645(.a(new_n838), .O(new_n839));
  nor2 g00646(.a(new_n808), .b(new_n802), .O(new_n840));
  nor2 g00647(.a(new_n840), .b(new_n839), .O(new_n841));
  inv1 g00648(.a(new_n840), .O(new_n842));
  nor2 g00649(.a(new_n842), .b(new_n838), .O(new_n843));
  nor2 g00650(.a(new_n843), .b(new_n841), .O(new_n844));
  inv1 g00651(.a(new_n844), .O(new_n845));
  nor2 g00652(.a(new_n438), .b(new_n257), .O(new_n846));
  inv1 g00653(.a(\a[16] ), .O(new_n847));
  nor2 g00654(.a(new_n847), .b(new_n198), .O(new_n848));
  nor2 g00655(.a(new_n848), .b(new_n846), .O(new_n849));
  nor2 g00656(.a(new_n847), .b(new_n257), .O(new_n850));
  inv1 g00657(.a(new_n850), .O(new_n851));
  nor2 g00658(.a(new_n851), .b(new_n442), .O(new_n852));
  nor2 g00659(.a(new_n852), .b(new_n849), .O(new_n853));
  nor2 g00660(.a(new_n853), .b(new_n541), .O(new_n854));
  inv1 g00661(.a(new_n853), .O(new_n855));
  nor2 g00662(.a(new_n855), .b(new_n540), .O(new_n856));
  nor2 g00663(.a(new_n856), .b(new_n854), .O(new_n857));
  nor2 g00664(.a(new_n857), .b(new_n845), .O(new_n858));
  inv1 g00665(.a(new_n857), .O(new_n859));
  nor2 g00666(.a(new_n859), .b(new_n844), .O(new_n860));
  nor2 g00667(.a(new_n860), .b(new_n858), .O(new_n861));
  nor2 g00668(.a(new_n861), .b(new_n837), .O(new_n862));
  inv1 g00669(.a(new_n861), .O(new_n863));
  nor2 g00670(.a(new_n863), .b(new_n836), .O(new_n864));
  nor2 g00671(.a(new_n864), .b(new_n862), .O(new_n865));
  inv1 g00672(.a(new_n773), .O(new_n866));
  nor2 g00673(.a(new_n363), .b(new_n295), .O(new_n867));
  nor2 g00674(.a(new_n800), .b(new_n194), .O(new_n868));
  nor2 g00675(.a(new_n868), .b(new_n867), .O(new_n869));
  inv1 g00676(.a(new_n867), .O(new_n870));
  inv1 g00677(.a(new_n868), .O(new_n871));
  nor2 g00678(.a(new_n871), .b(new_n870), .O(new_n872));
  nor2 g00679(.a(new_n872), .b(new_n869), .O(new_n873));
  inv1 g00680(.a(new_n873), .O(new_n874));
  nor2 g00681(.a(new_n874), .b(new_n866), .O(new_n875));
  nor2 g00682(.a(new_n873), .b(new_n773), .O(new_n876));
  nor2 g00683(.a(new_n876), .b(new_n875), .O(new_n877));
  inv1 g00684(.a(new_n877), .O(new_n878));
  nor2 g00685(.a(new_n762), .b(new_n755), .O(new_n879));
  inv1 g00686(.a(new_n879), .O(new_n880));
  nor2 g00687(.a(new_n880), .b(new_n878), .O(new_n881));
  nor2 g00688(.a(new_n879), .b(new_n877), .O(new_n882));
  nor2 g00689(.a(new_n882), .b(new_n881), .O(new_n883));
  inv1 g00690(.a(new_n883), .O(new_n884));
  nor2 g00691(.a(new_n569), .b(new_n214), .O(new_n885));
  inv1 g00692(.a(new_n885), .O(new_n886));
  nor2 g00693(.a(new_n613), .b(new_n203), .O(new_n887));
  nor2 g00694(.a(new_n699), .b(new_n196), .O(new_n888));
  nor2 g00695(.a(new_n888), .b(new_n887), .O(new_n889));
  nor2 g00696(.a(new_n699), .b(new_n203), .O(new_n890));
  inv1 g00697(.a(new_n890), .O(new_n891));
  nor2 g00698(.a(new_n891), .b(new_n752), .O(new_n892));
  nor2 g00699(.a(new_n892), .b(new_n889), .O(new_n893));
  nor2 g00700(.a(new_n893), .b(new_n886), .O(new_n894));
  inv1 g00701(.a(new_n893), .O(new_n895));
  nor2 g00702(.a(new_n895), .b(new_n885), .O(new_n896));
  nor2 g00703(.a(new_n896), .b(new_n894), .O(new_n897));
  nor2 g00704(.a(new_n811), .b(new_n794), .O(new_n898));
  inv1 g00705(.a(new_n898), .O(new_n899));
  nor2 g00706(.a(new_n899), .b(new_n897), .O(new_n900));
  inv1 g00707(.a(new_n897), .O(new_n901));
  nor2 g00708(.a(new_n898), .b(new_n901), .O(new_n902));
  nor2 g00709(.a(new_n902), .b(new_n900), .O(new_n903));
  inv1 g00710(.a(new_n903), .O(new_n904));
  nor2 g00711(.a(new_n904), .b(new_n884), .O(new_n905));
  nor2 g00712(.a(new_n903), .b(new_n883), .O(new_n906));
  nor2 g00713(.a(new_n906), .b(new_n905), .O(new_n907));
  nor2 g00714(.a(new_n907), .b(new_n865), .O(new_n908));
  inv1 g00715(.a(new_n865), .O(new_n909));
  inv1 g00716(.a(new_n907), .O(new_n910));
  nor2 g00717(.a(new_n910), .b(new_n909), .O(new_n911));
  nor2 g00718(.a(new_n911), .b(new_n908), .O(new_n912));
  inv1 g00719(.a(new_n912), .O(new_n913));
  nor2 g00720(.a(new_n913), .b(new_n835), .O(new_n914));
  inv1 g00721(.a(new_n835), .O(new_n915));
  nor2 g00722(.a(new_n912), .b(new_n915), .O(new_n916));
  nor2 g00723(.a(new_n916), .b(new_n914), .O(new_n917));
  nor2 g00724(.a(new_n830), .b(new_n825), .O(new_n918));
  inv1 g00725(.a(new_n918), .O(new_n919));
  nor2 g00726(.a(new_n919), .b(new_n917), .O(new_n920));
  inv1 g00727(.a(new_n917), .O(new_n921));
  nor2 g00728(.a(new_n918), .b(new_n921), .O(new_n922));
  nor2 g00729(.a(new_n922), .b(new_n920), .O(new_n923));
  inv1 g00730(.a(new_n923), .O(\asquared[17] ));
  nor2 g00731(.a(new_n911), .b(new_n864), .O(new_n925));
  nor2 g00732(.a(new_n905), .b(new_n900), .O(new_n926));
  inv1 g00733(.a(new_n926), .O(new_n927));
  nor2 g00734(.a(new_n363), .b(new_n322), .O(new_n928));
  nor2 g00735(.a(new_n438), .b(new_n295), .O(new_n929));
  nor2 g00736(.a(new_n929), .b(new_n928), .O(new_n930));
  nor2 g00737(.a(new_n438), .b(new_n322), .O(new_n931));
  inv1 g00738(.a(new_n931), .O(new_n932));
  nor2 g00739(.a(new_n932), .b(new_n870), .O(new_n933));
  nor2 g00740(.a(new_n933), .b(new_n930), .O(new_n934));
  nor2 g00741(.a(new_n934), .b(new_n891), .O(new_n935));
  inv1 g00742(.a(new_n934), .O(new_n936));
  nor2 g00743(.a(new_n936), .b(new_n890), .O(new_n937));
  nor2 g00744(.a(new_n937), .b(new_n935), .O(new_n938));
  inv1 g00745(.a(new_n872), .O(new_n939));
  nor2 g00746(.a(new_n569), .b(new_n229), .O(new_n940));
  inv1 g00747(.a(\a[17] ), .O(new_n941));
  nor2 g00748(.a(new_n941), .b(new_n198), .O(new_n942));
  nor2 g00749(.a(new_n942), .b(new_n940), .O(new_n943));
  inv1 g00750(.a(new_n940), .O(new_n944));
  inv1 g00751(.a(new_n942), .O(new_n945));
  nor2 g00752(.a(new_n945), .b(new_n944), .O(new_n946));
  nor2 g00753(.a(new_n946), .b(new_n943), .O(new_n947));
  inv1 g00754(.a(new_n947), .O(new_n948));
  nor2 g00755(.a(new_n948), .b(new_n939), .O(new_n949));
  nor2 g00756(.a(new_n947), .b(new_n872), .O(new_n950));
  nor2 g00757(.a(new_n950), .b(new_n949), .O(new_n951));
  inv1 g00758(.a(new_n951), .O(new_n952));
  nor2 g00759(.a(new_n952), .b(new_n938), .O(new_n953));
  inv1 g00760(.a(new_n938), .O(new_n954));
  nor2 g00761(.a(new_n951), .b(new_n954), .O(new_n955));
  nor2 g00762(.a(new_n955), .b(new_n953), .O(new_n956));
  inv1 g00763(.a(new_n956), .O(new_n957));
  nor2 g00764(.a(new_n502), .b(new_n257), .O(new_n958));
  inv1 g00765(.a(new_n958), .O(new_n959));
  nor2 g00766(.a(new_n800), .b(new_n196), .O(new_n960));
  nor2 g00767(.a(new_n960), .b(new_n616), .O(new_n961));
  nor2 g00768(.a(new_n800), .b(new_n214), .O(new_n962));
  inv1 g00769(.a(new_n962), .O(new_n963));
  nor2 g00770(.a(new_n963), .b(new_n752), .O(new_n964));
  nor2 g00771(.a(new_n964), .b(new_n961), .O(new_n965));
  nor2 g00772(.a(new_n965), .b(new_n959), .O(new_n966));
  inv1 g00773(.a(new_n965), .O(new_n967));
  nor2 g00774(.a(new_n967), .b(new_n958), .O(new_n968));
  nor2 g00775(.a(new_n968), .b(new_n966), .O(new_n969));
  nor2 g00776(.a(new_n969), .b(new_n957), .O(new_n970));
  inv1 g00777(.a(new_n969), .O(new_n971));
  nor2 g00778(.a(new_n971), .b(new_n956), .O(new_n972));
  nor2 g00779(.a(new_n972), .b(new_n970), .O(new_n973));
  nor2 g00780(.a(new_n973), .b(new_n927), .O(new_n974));
  inv1 g00781(.a(new_n973), .O(new_n975));
  nor2 g00782(.a(new_n975), .b(new_n926), .O(new_n976));
  nor2 g00783(.a(new_n976), .b(new_n974), .O(new_n977));
  inv1 g00784(.a(new_n977), .O(new_n978));
  nor2 g00785(.a(new_n881), .b(new_n875), .O(new_n979));
  inv1 g00786(.a(new_n979), .O(new_n980));
  nor2 g00787(.a(new_n858), .b(new_n843), .O(new_n981));
  inv1 g00788(.a(new_n981), .O(new_n982));
  nor2 g00789(.a(new_n982), .b(new_n980), .O(new_n983));
  nor2 g00790(.a(new_n981), .b(new_n979), .O(new_n984));
  nor2 g00791(.a(new_n984), .b(new_n983), .O(new_n985));
  nor2 g00792(.a(new_n847), .b(new_n194), .O(new_n986));
  nor2 g00793(.a(new_n986), .b(\a[9] ), .O(new_n987));
  nor2 g00794(.a(new_n847), .b(new_n363), .O(new_n988));
  inv1 g00795(.a(new_n988), .O(new_n989));
  nor2 g00796(.a(new_n989), .b(new_n194), .O(new_n990));
  nor2 g00797(.a(new_n990), .b(new_n987), .O(new_n991));
  inv1 g00798(.a(new_n991), .O(new_n992));
  nor2 g00799(.a(new_n896), .b(new_n889), .O(new_n993));
  inv1 g00800(.a(new_n993), .O(new_n994));
  nor2 g00801(.a(new_n994), .b(new_n992), .O(new_n995));
  nor2 g00802(.a(new_n993), .b(new_n991), .O(new_n996));
  nor2 g00803(.a(new_n996), .b(new_n995), .O(new_n997));
  inv1 g00804(.a(new_n997), .O(new_n998));
  nor2 g00805(.a(new_n856), .b(new_n849), .O(new_n999));
  inv1 g00806(.a(new_n999), .O(new_n1000));
  nor2 g00807(.a(new_n1000), .b(new_n998), .O(new_n1001));
  nor2 g00808(.a(new_n999), .b(new_n997), .O(new_n1002));
  nor2 g00809(.a(new_n1002), .b(new_n1001), .O(new_n1003));
  nor2 g00810(.a(new_n1003), .b(new_n985), .O(new_n1004));
  inv1 g00811(.a(new_n985), .O(new_n1005));
  inv1 g00812(.a(new_n1003), .O(new_n1006));
  nor2 g00813(.a(new_n1006), .b(new_n1005), .O(new_n1007));
  nor2 g00814(.a(new_n1007), .b(new_n1004), .O(new_n1008));
  inv1 g00815(.a(new_n1008), .O(new_n1009));
  nor2 g00816(.a(new_n1009), .b(new_n978), .O(new_n1010));
  nor2 g00817(.a(new_n1008), .b(new_n977), .O(new_n1011));
  nor2 g00818(.a(new_n1011), .b(new_n1010), .O(new_n1012));
  inv1 g00819(.a(new_n1012), .O(new_n1013));
  nor2 g00820(.a(new_n1013), .b(new_n925), .O(new_n1014));
  inv1 g00821(.a(new_n925), .O(new_n1015));
  nor2 g00822(.a(new_n1012), .b(new_n1015), .O(new_n1016));
  nor2 g00823(.a(new_n1016), .b(new_n1014), .O(new_n1017));
  inv1 g00824(.a(new_n1017), .O(new_n1018));
  nor2 g00825(.a(new_n918), .b(new_n914), .O(new_n1019));
  nor2 g00826(.a(new_n1019), .b(new_n916), .O(new_n1020));
  inv1 g00827(.a(new_n1020), .O(new_n1021));
  nor2 g00828(.a(new_n1021), .b(new_n1018), .O(new_n1022));
  nor2 g00829(.a(new_n1020), .b(new_n1017), .O(new_n1023));
  nor2 g00830(.a(new_n1023), .b(new_n1022), .O(\asquared[18] ));
  nor2 g00831(.a(new_n1010), .b(new_n976), .O(new_n1025));
  nor2 g00832(.a(new_n949), .b(new_n946), .O(new_n1026));
  inv1 g00833(.a(new_n1026), .O(new_n1027));
  nor2 g00834(.a(new_n937), .b(new_n930), .O(new_n1028));
  nor2 g00835(.a(new_n968), .b(new_n961), .O(new_n1029));
  nor2 g00836(.a(new_n1029), .b(new_n1028), .O(new_n1030));
  inv1 g00837(.a(new_n1028), .O(new_n1031));
  inv1 g00838(.a(new_n1029), .O(new_n1032));
  nor2 g00839(.a(new_n1032), .b(new_n1031), .O(new_n1033));
  nor2 g00840(.a(new_n1033), .b(new_n1030), .O(new_n1034));
  nor2 g00841(.a(new_n1034), .b(new_n1027), .O(new_n1035));
  inv1 g00842(.a(new_n1034), .O(new_n1036));
  nor2 g00843(.a(new_n1036), .b(new_n1026), .O(new_n1037));
  nor2 g00844(.a(new_n1037), .b(new_n1035), .O(new_n1038));
  inv1 g00845(.a(new_n1038), .O(new_n1039));
  nor2 g00846(.a(new_n1001), .b(new_n995), .O(new_n1040));
  inv1 g00847(.a(new_n1040), .O(new_n1041));
  nor2 g00848(.a(new_n970), .b(new_n953), .O(new_n1042));
  inv1 g00849(.a(new_n1042), .O(new_n1043));
  nor2 g00850(.a(new_n1043), .b(new_n1041), .O(new_n1044));
  nor2 g00851(.a(new_n1042), .b(new_n1040), .O(new_n1045));
  nor2 g00852(.a(new_n1045), .b(new_n1044), .O(new_n1046));
  inv1 g00853(.a(new_n1046), .O(new_n1047));
  nor2 g00854(.a(new_n1047), .b(new_n1039), .O(new_n1048));
  nor2 g00855(.a(new_n1046), .b(new_n1038), .O(new_n1049));
  nor2 g00856(.a(new_n1049), .b(new_n1048), .O(new_n1050));
  inv1 g00857(.a(new_n1050), .O(new_n1051));
  nor2 g00858(.a(new_n1007), .b(new_n984), .O(new_n1052));
  nor2 g00859(.a(new_n569), .b(new_n257), .O(new_n1053));
  nor2 g00860(.a(new_n1053), .b(new_n990), .O(new_n1054));
  inv1 g00861(.a(new_n990), .O(new_n1055));
  inv1 g00862(.a(new_n1053), .O(new_n1056));
  nor2 g00863(.a(new_n1056), .b(new_n1055), .O(new_n1057));
  nor2 g00864(.a(new_n1057), .b(new_n1054), .O(new_n1058));
  inv1 g00865(.a(new_n1058), .O(new_n1059));
  nor2 g00866(.a(new_n941), .b(new_n194), .O(new_n1060));
  inv1 g00867(.a(new_n1060), .O(new_n1061));
  nor2 g00868(.a(new_n1061), .b(new_n932), .O(new_n1062));
  nor2 g00869(.a(new_n1060), .b(new_n931), .O(new_n1063));
  nor2 g00870(.a(new_n1063), .b(new_n1062), .O(new_n1064));
  inv1 g00871(.a(new_n1064), .O(new_n1065));
  nor2 g00872(.a(new_n1065), .b(new_n1059), .O(new_n1066));
  nor2 g00873(.a(new_n1064), .b(new_n1058), .O(new_n1067));
  nor2 g00874(.a(new_n1067), .b(new_n1066), .O(new_n1068));
  inv1 g00875(.a(new_n1068), .O(new_n1069));
  nor2 g00876(.a(new_n699), .b(new_n214), .O(new_n1070));
  inv1 g00877(.a(new_n1070), .O(new_n1071));
  nor2 g00878(.a(new_n800), .b(new_n203), .O(new_n1072));
  nor2 g00879(.a(new_n847), .b(new_n196), .O(new_n1073));
  nor2 g00880(.a(new_n1073), .b(new_n1072), .O(new_n1074));
  inv1 g00881(.a(new_n960), .O(new_n1075));
  nor2 g00882(.a(new_n847), .b(new_n203), .O(new_n1076));
  inv1 g00883(.a(new_n1076), .O(new_n1077));
  nor2 g00884(.a(new_n1077), .b(new_n1075), .O(new_n1078));
  nor2 g00885(.a(new_n1078), .b(new_n1074), .O(new_n1079));
  nor2 g00886(.a(new_n1079), .b(new_n1071), .O(new_n1080));
  inv1 g00887(.a(new_n1079), .O(new_n1081));
  nor2 g00888(.a(new_n1081), .b(new_n1070), .O(new_n1082));
  nor2 g00889(.a(new_n1082), .b(new_n1080), .O(new_n1083));
  nor2 g00890(.a(new_n502), .b(new_n295), .O(new_n1084));
  inv1 g00891(.a(new_n1084), .O(new_n1085));
  inv1 g00892(.a(\a[18] ), .O(new_n1086));
  nor2 g00893(.a(new_n1086), .b(new_n198), .O(new_n1087));
  nor2 g00894(.a(new_n613), .b(new_n229), .O(new_n1088));
  nor2 g00895(.a(new_n1088), .b(new_n1087), .O(new_n1089));
  inv1 g00896(.a(new_n1087), .O(new_n1090));
  inv1 g00897(.a(new_n1088), .O(new_n1091));
  nor2 g00898(.a(new_n1091), .b(new_n1090), .O(new_n1092));
  nor2 g00899(.a(new_n1092), .b(new_n1089), .O(new_n1093));
  nor2 g00900(.a(new_n1093), .b(new_n1085), .O(new_n1094));
  inv1 g00901(.a(new_n1093), .O(new_n1095));
  nor2 g00902(.a(new_n1095), .b(new_n1084), .O(new_n1096));
  nor2 g00903(.a(new_n1096), .b(new_n1094), .O(new_n1097));
  nor2 g00904(.a(new_n1097), .b(new_n1083), .O(new_n1098));
  inv1 g00905(.a(new_n1083), .O(new_n1099));
  inv1 g00906(.a(new_n1097), .O(new_n1100));
  nor2 g00907(.a(new_n1100), .b(new_n1099), .O(new_n1101));
  nor2 g00908(.a(new_n1101), .b(new_n1098), .O(new_n1102));
  inv1 g00909(.a(new_n1102), .O(new_n1103));
  nor2 g00910(.a(new_n1103), .b(new_n1069), .O(new_n1104));
  nor2 g00911(.a(new_n1102), .b(new_n1068), .O(new_n1105));
  nor2 g00912(.a(new_n1105), .b(new_n1104), .O(new_n1106));
  inv1 g00913(.a(new_n1106), .O(new_n1107));
  nor2 g00914(.a(new_n1107), .b(new_n1052), .O(new_n1108));
  inv1 g00915(.a(new_n1052), .O(new_n1109));
  nor2 g00916(.a(new_n1106), .b(new_n1109), .O(new_n1110));
  nor2 g00917(.a(new_n1110), .b(new_n1108), .O(new_n1111));
  inv1 g00918(.a(new_n1111), .O(new_n1112));
  nor2 g00919(.a(new_n1112), .b(new_n1051), .O(new_n1113));
  nor2 g00920(.a(new_n1111), .b(new_n1050), .O(new_n1114));
  nor2 g00921(.a(new_n1114), .b(new_n1113), .O(new_n1115));
  inv1 g00922(.a(new_n1115), .O(new_n1116));
  nor2 g00923(.a(new_n1116), .b(new_n1025), .O(new_n1117));
  inv1 g00924(.a(new_n1025), .O(new_n1118));
  nor2 g00925(.a(new_n1115), .b(new_n1118), .O(new_n1119));
  nor2 g00926(.a(new_n1119), .b(new_n1117), .O(new_n1120));
  inv1 g00927(.a(new_n1120), .O(new_n1121));
  nor2 g00928(.a(new_n1020), .b(new_n1014), .O(new_n1122));
  nor2 g00929(.a(new_n1122), .b(new_n1016), .O(new_n1123));
  inv1 g00930(.a(new_n1123), .O(new_n1124));
  nor2 g00931(.a(new_n1124), .b(new_n1121), .O(new_n1125));
  nor2 g00932(.a(new_n1123), .b(new_n1120), .O(new_n1126));
  nor2 g00933(.a(new_n1126), .b(new_n1125), .O(\asquared[19] ));
  nor2 g00934(.a(new_n1104), .b(new_n1098), .O(new_n1128));
  nor2 g00935(.a(new_n1086), .b(new_n194), .O(new_n1129));
  nor2 g00936(.a(new_n1129), .b(\a[10] ), .O(new_n1130));
  inv1 g00937(.a(new_n1129), .O(new_n1131));
  nor2 g00938(.a(new_n1131), .b(new_n438), .O(new_n1132));
  nor2 g00939(.a(new_n1132), .b(new_n1130), .O(new_n1133));
  nor2 g00940(.a(new_n1133), .b(new_n1062), .O(new_n1134));
  inv1 g00941(.a(new_n1062), .O(new_n1135));
  nor2 g00942(.a(new_n1135), .b(\a[18] ), .O(new_n1136));
  nor2 g00943(.a(new_n1136), .b(new_n1134), .O(new_n1137));
  inv1 g00944(.a(new_n1137), .O(new_n1138));
  nor2 g00945(.a(new_n1082), .b(new_n1074), .O(new_n1139));
  inv1 g00946(.a(new_n1139), .O(new_n1140));
  nor2 g00947(.a(new_n1140), .b(new_n1138), .O(new_n1141));
  nor2 g00948(.a(new_n1139), .b(new_n1137), .O(new_n1142));
  nor2 g00949(.a(new_n1142), .b(new_n1141), .O(new_n1143));
  inv1 g00950(.a(new_n1143), .O(new_n1144));
  nor2 g00951(.a(new_n1144), .b(new_n1128), .O(new_n1145));
  inv1 g00952(.a(new_n1128), .O(new_n1146));
  nor2 g00953(.a(new_n1143), .b(new_n1146), .O(new_n1147));
  nor2 g00954(.a(new_n1147), .b(new_n1145), .O(new_n1148));
  inv1 g00955(.a(new_n1148), .O(new_n1149));
  nor2 g00956(.a(new_n1066), .b(new_n1057), .O(new_n1150));
  inv1 g00957(.a(new_n1150), .O(new_n1151));
  nor2 g00958(.a(new_n1096), .b(new_n1089), .O(new_n1152));
  nor2 g00959(.a(new_n1152), .b(new_n1151), .O(new_n1153));
  inv1 g00960(.a(new_n1152), .O(new_n1154));
  nor2 g00961(.a(new_n1154), .b(new_n1150), .O(new_n1155));
  nor2 g00962(.a(new_n1155), .b(new_n1153), .O(new_n1156));
  inv1 g00963(.a(new_n1156), .O(new_n1157));
  nor2 g00964(.a(new_n438), .b(new_n363), .O(new_n1158));
  nor2 g00965(.a(new_n502), .b(new_n322), .O(new_n1159));
  nor2 g00966(.a(new_n1159), .b(new_n1158), .O(new_n1160));
  inv1 g00967(.a(new_n1158), .O(new_n1161));
  inv1 g00968(.a(new_n1159), .O(new_n1162));
  nor2 g00969(.a(new_n1162), .b(new_n1161), .O(new_n1163));
  nor2 g00970(.a(new_n1163), .b(new_n1160), .O(new_n1164));
  nor2 g00971(.a(new_n1164), .b(new_n1077), .O(new_n1165));
  inv1 g00972(.a(new_n1164), .O(new_n1166));
  nor2 g00973(.a(new_n1166), .b(new_n1076), .O(new_n1167));
  nor2 g00974(.a(new_n1167), .b(new_n1165), .O(new_n1168));
  nor2 g00975(.a(new_n1168), .b(new_n1157), .O(new_n1169));
  inv1 g00976(.a(new_n1168), .O(new_n1170));
  nor2 g00977(.a(new_n1170), .b(new_n1156), .O(new_n1171));
  nor2 g00978(.a(new_n1171), .b(new_n1169), .O(new_n1172));
  inv1 g00979(.a(new_n1172), .O(new_n1173));
  nor2 g00980(.a(new_n1173), .b(new_n1149), .O(new_n1174));
  nor2 g00981(.a(new_n1172), .b(new_n1148), .O(new_n1175));
  nor2 g00982(.a(new_n1175), .b(new_n1174), .O(new_n1176));
  inv1 g00983(.a(new_n1176), .O(new_n1177));
  nor2 g00984(.a(new_n1037), .b(new_n1033), .O(new_n1178));
  inv1 g00985(.a(new_n1178), .O(new_n1179));
  nor2 g00986(.a(new_n699), .b(new_n229), .O(new_n1180));
  inv1 g00987(.a(new_n1180), .O(new_n1181));
  nor2 g00988(.a(new_n613), .b(new_n257), .O(new_n1182));
  nor2 g00989(.a(new_n569), .b(new_n295), .O(new_n1183));
  nor2 g00990(.a(new_n1183), .b(new_n1182), .O(new_n1184));
  nor2 g00991(.a(new_n613), .b(new_n295), .O(new_n1185));
  inv1 g00992(.a(new_n1185), .O(new_n1186));
  nor2 g00993(.a(new_n1186), .b(new_n1056), .O(new_n1187));
  nor2 g00994(.a(new_n1187), .b(new_n1184), .O(new_n1188));
  nor2 g00995(.a(new_n1188), .b(new_n1181), .O(new_n1189));
  inv1 g00996(.a(new_n1188), .O(new_n1190));
  nor2 g00997(.a(new_n1190), .b(new_n1180), .O(new_n1191));
  nor2 g00998(.a(new_n1191), .b(new_n1189), .O(new_n1192));
  nor2 g00999(.a(new_n941), .b(new_n196), .O(new_n1193));
  nor2 g01000(.a(new_n1193), .b(new_n962), .O(new_n1194));
  nor2 g01001(.a(new_n941), .b(new_n214), .O(new_n1195));
  inv1 g01002(.a(new_n1195), .O(new_n1196));
  nor2 g01003(.a(new_n1196), .b(new_n1075), .O(new_n1197));
  nor2 g01004(.a(new_n1197), .b(new_n1194), .O(new_n1198));
  inv1 g01005(.a(\a[19] ), .O(new_n1199));
  nor2 g01006(.a(new_n1199), .b(new_n198), .O(new_n1200));
  inv1 g01007(.a(new_n1200), .O(new_n1201));
  nor2 g01008(.a(new_n1201), .b(new_n1198), .O(new_n1202));
  inv1 g01009(.a(new_n1198), .O(new_n1203));
  nor2 g01010(.a(new_n1200), .b(new_n1203), .O(new_n1204));
  nor2 g01011(.a(new_n1204), .b(new_n1202), .O(new_n1205));
  nor2 g01012(.a(new_n1205), .b(new_n1192), .O(new_n1206));
  inv1 g01013(.a(new_n1192), .O(new_n1207));
  inv1 g01014(.a(new_n1205), .O(new_n1208));
  nor2 g01015(.a(new_n1208), .b(new_n1207), .O(new_n1209));
  nor2 g01016(.a(new_n1209), .b(new_n1206), .O(new_n1210));
  nor2 g01017(.a(new_n1210), .b(new_n1179), .O(new_n1211));
  inv1 g01018(.a(new_n1210), .O(new_n1212));
  nor2 g01019(.a(new_n1212), .b(new_n1178), .O(new_n1213));
  nor2 g01020(.a(new_n1213), .b(new_n1211), .O(new_n1214));
  inv1 g01021(.a(new_n1214), .O(new_n1215));
  nor2 g01022(.a(new_n1048), .b(new_n1045), .O(new_n1216));
  nor2 g01023(.a(new_n1216), .b(new_n1215), .O(new_n1217));
  inv1 g01024(.a(new_n1216), .O(new_n1218));
  nor2 g01025(.a(new_n1218), .b(new_n1214), .O(new_n1219));
  nor2 g01026(.a(new_n1219), .b(new_n1217), .O(new_n1220));
  inv1 g01027(.a(new_n1220), .O(new_n1221));
  nor2 g01028(.a(new_n1221), .b(new_n1177), .O(new_n1222));
  nor2 g01029(.a(new_n1220), .b(new_n1176), .O(new_n1223));
  nor2 g01030(.a(new_n1223), .b(new_n1222), .O(new_n1224));
  nor2 g01031(.a(new_n1113), .b(new_n1108), .O(new_n1225));
  inv1 g01032(.a(new_n1225), .O(new_n1226));
  nor2 g01033(.a(new_n1226), .b(new_n1224), .O(new_n1227));
  inv1 g01034(.a(new_n1224), .O(new_n1228));
  nor2 g01035(.a(new_n1225), .b(new_n1228), .O(new_n1229));
  nor2 g01036(.a(new_n1229), .b(new_n1227), .O(new_n1230));
  inv1 g01037(.a(new_n1230), .O(new_n1231));
  nor2 g01038(.a(new_n1123), .b(new_n1117), .O(new_n1232));
  nor2 g01039(.a(new_n1232), .b(new_n1119), .O(new_n1233));
  nor2 g01040(.a(new_n1233), .b(new_n1231), .O(new_n1234));
  inv1 g01041(.a(new_n1233), .O(new_n1235));
  nor2 g01042(.a(new_n1235), .b(new_n1230), .O(new_n1236));
  nor2 g01043(.a(new_n1236), .b(new_n1234), .O(new_n1237));
  inv1 g01044(.a(new_n1237), .O(\asquared[20] ));
  nor2 g01045(.a(new_n1222), .b(new_n1217), .O(new_n1239));
  nor2 g01046(.a(new_n1141), .b(new_n1136), .O(new_n1240));
  nor2 g01047(.a(new_n1086), .b(new_n196), .O(new_n1241));
  inv1 g01048(.a(new_n1241), .O(new_n1242));
  nor2 g01049(.a(new_n941), .b(new_n203), .O(new_n1243));
  nor2 g01050(.a(new_n847), .b(new_n214), .O(new_n1244));
  nor2 g01051(.a(new_n1244), .b(new_n1243), .O(new_n1245));
  nor2 g01052(.a(new_n1196), .b(new_n1077), .O(new_n1246));
  nor2 g01053(.a(new_n1246), .b(new_n1245), .O(new_n1247));
  nor2 g01054(.a(new_n1247), .b(new_n1242), .O(new_n1248));
  inv1 g01055(.a(new_n1247), .O(new_n1249));
  nor2 g01056(.a(new_n1249), .b(new_n1241), .O(new_n1250));
  nor2 g01057(.a(new_n1250), .b(new_n1248), .O(new_n1251));
  nor2 g01058(.a(new_n1251), .b(new_n1240), .O(new_n1252));
  inv1 g01059(.a(new_n1240), .O(new_n1253));
  inv1 g01060(.a(new_n1251), .O(new_n1254));
  nor2 g01061(.a(new_n1254), .b(new_n1253), .O(new_n1255));
  nor2 g01062(.a(new_n1255), .b(new_n1252), .O(new_n1256));
  nor2 g01063(.a(new_n1169), .b(new_n1155), .O(new_n1257));
  inv1 g01064(.a(new_n1257), .O(new_n1258));
  nor2 g01065(.a(new_n1258), .b(new_n1256), .O(new_n1259));
  inv1 g01066(.a(new_n1256), .O(new_n1260));
  nor2 g01067(.a(new_n1257), .b(new_n1260), .O(new_n1261));
  nor2 g01068(.a(new_n1261), .b(new_n1259), .O(new_n1262));
  nor2 g01069(.a(new_n1174), .b(new_n1145), .O(new_n1263));
  inv1 g01070(.a(new_n1263), .O(new_n1264));
  nor2 g01071(.a(new_n1264), .b(new_n1262), .O(new_n1265));
  inv1 g01072(.a(new_n1262), .O(new_n1266));
  nor2 g01073(.a(new_n1263), .b(new_n1266), .O(new_n1267));
  nor2 g01074(.a(new_n1267), .b(new_n1265), .O(new_n1268));
  inv1 g01075(.a(new_n1268), .O(new_n1269));
  nor2 g01076(.a(new_n1213), .b(new_n1206), .O(new_n1270));
  inv1 g01077(.a(new_n1270), .O(new_n1271));
  nor2 g01078(.a(new_n502), .b(new_n363), .O(new_n1272));
  nor2 g01079(.a(new_n1199), .b(new_n194), .O(new_n1273));
  nor2 g01080(.a(new_n1273), .b(new_n1272), .O(new_n1274));
  inv1 g01081(.a(new_n1272), .O(new_n1275));
  inv1 g01082(.a(new_n1273), .O(new_n1276));
  nor2 g01083(.a(new_n1276), .b(new_n1275), .O(new_n1277));
  nor2 g01084(.a(new_n1277), .b(new_n1274), .O(new_n1278));
  inv1 g01085(.a(new_n1278), .O(new_n1279));
  nor2 g01086(.a(new_n1167), .b(new_n1160), .O(new_n1280));
  inv1 g01087(.a(new_n1280), .O(new_n1281));
  nor2 g01088(.a(new_n1281), .b(new_n1279), .O(new_n1282));
  nor2 g01089(.a(new_n1280), .b(new_n1278), .O(new_n1283));
  nor2 g01090(.a(new_n1283), .b(new_n1282), .O(new_n1284));
  inv1 g01091(.a(new_n1284), .O(new_n1285));
  nor2 g01092(.a(new_n1204), .b(new_n1194), .O(new_n1286));
  inv1 g01093(.a(new_n1286), .O(new_n1287));
  nor2 g01094(.a(new_n1287), .b(new_n1285), .O(new_n1288));
  nor2 g01095(.a(new_n1286), .b(new_n1284), .O(new_n1289));
  nor2 g01096(.a(new_n1289), .b(new_n1288), .O(new_n1290));
  nor2 g01097(.a(new_n1290), .b(new_n1271), .O(new_n1291));
  inv1 g01098(.a(new_n1290), .O(new_n1292));
  nor2 g01099(.a(new_n1292), .b(new_n1270), .O(new_n1293));
  nor2 g01100(.a(new_n1293), .b(new_n1291), .O(new_n1294));
  inv1 g01101(.a(new_n1294), .O(new_n1295));
  inv1 g01102(.a(new_n1132), .O(new_n1296));
  inv1 g01103(.a(\a[20] ), .O(new_n1297));
  nor2 g01104(.a(new_n1297), .b(new_n198), .O(new_n1298));
  nor2 g01105(.a(new_n1298), .b(new_n1185), .O(new_n1299));
  inv1 g01106(.a(new_n1298), .O(new_n1300));
  nor2 g01107(.a(new_n1300), .b(new_n1186), .O(new_n1301));
  nor2 g01108(.a(new_n1301), .b(new_n1299), .O(new_n1302));
  inv1 g01109(.a(new_n1302), .O(new_n1303));
  nor2 g01110(.a(new_n1303), .b(new_n1296), .O(new_n1304));
  nor2 g01111(.a(new_n1302), .b(new_n1132), .O(new_n1305));
  nor2 g01112(.a(new_n1305), .b(new_n1304), .O(new_n1306));
  inv1 g01113(.a(new_n1306), .O(new_n1307));
  nor2 g01114(.a(new_n1191), .b(new_n1184), .O(new_n1308));
  inv1 g01115(.a(new_n1308), .O(new_n1309));
  nor2 g01116(.a(new_n1309), .b(new_n1307), .O(new_n1310));
  nor2 g01117(.a(new_n1308), .b(new_n1306), .O(new_n1311));
  nor2 g01118(.a(new_n1311), .b(new_n1310), .O(new_n1312));
  inv1 g01119(.a(new_n1312), .O(new_n1313));
  nor2 g01120(.a(new_n569), .b(new_n322), .O(new_n1314));
  inv1 g01121(.a(new_n1314), .O(new_n1315));
  nor2 g01122(.a(new_n800), .b(new_n229), .O(new_n1316));
  nor2 g01123(.a(new_n699), .b(new_n257), .O(new_n1317));
  nor2 g01124(.a(new_n1317), .b(new_n1316), .O(new_n1318));
  nor2 g01125(.a(new_n800), .b(new_n257), .O(new_n1319));
  inv1 g01126(.a(new_n1319), .O(new_n1320));
  nor2 g01127(.a(new_n1320), .b(new_n1181), .O(new_n1321));
  nor2 g01128(.a(new_n1321), .b(new_n1318), .O(new_n1322));
  nor2 g01129(.a(new_n1322), .b(new_n1315), .O(new_n1323));
  inv1 g01130(.a(new_n1322), .O(new_n1324));
  nor2 g01131(.a(new_n1324), .b(new_n1314), .O(new_n1325));
  nor2 g01132(.a(new_n1325), .b(new_n1323), .O(new_n1326));
  nor2 g01133(.a(new_n1326), .b(new_n1313), .O(new_n1327));
  inv1 g01134(.a(new_n1326), .O(new_n1328));
  nor2 g01135(.a(new_n1328), .b(new_n1312), .O(new_n1329));
  nor2 g01136(.a(new_n1329), .b(new_n1327), .O(new_n1330));
  inv1 g01137(.a(new_n1330), .O(new_n1331));
  nor2 g01138(.a(new_n1331), .b(new_n1295), .O(new_n1332));
  nor2 g01139(.a(new_n1330), .b(new_n1294), .O(new_n1333));
  nor2 g01140(.a(new_n1333), .b(new_n1332), .O(new_n1334));
  inv1 g01141(.a(new_n1334), .O(new_n1335));
  nor2 g01142(.a(new_n1335), .b(new_n1269), .O(new_n1336));
  nor2 g01143(.a(new_n1334), .b(new_n1268), .O(new_n1337));
  nor2 g01144(.a(new_n1337), .b(new_n1336), .O(new_n1338));
  inv1 g01145(.a(new_n1338), .O(new_n1339));
  nor2 g01146(.a(new_n1339), .b(new_n1239), .O(new_n1340));
  inv1 g01147(.a(new_n1239), .O(new_n1341));
  nor2 g01148(.a(new_n1338), .b(new_n1341), .O(new_n1342));
  nor2 g01149(.a(new_n1342), .b(new_n1340), .O(new_n1343));
  inv1 g01150(.a(new_n1343), .O(new_n1344));
  nor2 g01151(.a(new_n1234), .b(new_n1227), .O(new_n1345));
  nor2 g01152(.a(new_n1345), .b(new_n1344), .O(new_n1346));
  inv1 g01153(.a(new_n1345), .O(new_n1347));
  nor2 g01154(.a(new_n1347), .b(new_n1343), .O(new_n1348));
  nor2 g01155(.a(new_n1348), .b(new_n1346), .O(new_n1349));
  inv1 g01156(.a(new_n1349), .O(\asquared[21] ));
  nor2 g01157(.a(new_n1336), .b(new_n1267), .O(new_n1351));
  nor2 g01158(.a(new_n1250), .b(new_n1245), .O(new_n1352));
  nor2 g01159(.a(new_n1325), .b(new_n1318), .O(new_n1353));
  nor2 g01160(.a(new_n1353), .b(new_n1352), .O(new_n1354));
  inv1 g01161(.a(new_n1352), .O(new_n1355));
  inv1 g01162(.a(new_n1353), .O(new_n1356));
  nor2 g01163(.a(new_n1356), .b(new_n1355), .O(new_n1357));
  nor2 g01164(.a(new_n1357), .b(new_n1354), .O(new_n1358));
  nor2 g01165(.a(new_n1304), .b(new_n1301), .O(new_n1359));
  inv1 g01166(.a(new_n1359), .O(new_n1360));
  nor2 g01167(.a(new_n1360), .b(new_n1358), .O(new_n1361));
  inv1 g01168(.a(new_n1358), .O(new_n1362));
  nor2 g01169(.a(new_n1359), .b(new_n1362), .O(new_n1363));
  nor2 g01170(.a(new_n1363), .b(new_n1361), .O(new_n1364));
  nor2 g01171(.a(new_n1261), .b(new_n1252), .O(new_n1365));
  inv1 g01172(.a(new_n1365), .O(new_n1366));
  nor2 g01173(.a(new_n1366), .b(new_n1364), .O(new_n1367));
  inv1 g01174(.a(new_n1364), .O(new_n1368));
  nor2 g01175(.a(new_n1365), .b(new_n1368), .O(new_n1369));
  nor2 g01176(.a(new_n1369), .b(new_n1367), .O(new_n1370));
  nor2 g01177(.a(new_n502), .b(new_n438), .O(new_n1371));
  nor2 g01178(.a(new_n569), .b(new_n363), .O(new_n1372));
  nor2 g01179(.a(new_n1372), .b(new_n1371), .O(new_n1373));
  nor2 g01180(.a(new_n569), .b(new_n438), .O(new_n1374));
  inv1 g01181(.a(new_n1374), .O(new_n1375));
  nor2 g01182(.a(new_n1375), .b(new_n1275), .O(new_n1376));
  nor2 g01183(.a(new_n1376), .b(new_n1373), .O(new_n1377));
  nor2 g01184(.a(new_n1377), .b(new_n1196), .O(new_n1378));
  inv1 g01185(.a(new_n1377), .O(new_n1379));
  nor2 g01186(.a(new_n1379), .b(new_n1195), .O(new_n1380));
  nor2 g01187(.a(new_n1380), .b(new_n1378), .O(new_n1381));
  inv1 g01188(.a(new_n1381), .O(new_n1382));
  nor2 g01189(.a(new_n613), .b(new_n322), .O(new_n1383));
  nor2 g01190(.a(new_n699), .b(new_n295), .O(new_n1384));
  nor2 g01191(.a(new_n1384), .b(new_n1383), .O(new_n1385));
  nor2 g01192(.a(new_n699), .b(new_n322), .O(new_n1386));
  inv1 g01193(.a(new_n1386), .O(new_n1387));
  nor2 g01194(.a(new_n1387), .b(new_n1186), .O(new_n1388));
  nor2 g01195(.a(new_n1388), .b(new_n1385), .O(new_n1389));
  nor2 g01196(.a(new_n1389), .b(new_n1320), .O(new_n1390));
  inv1 g01197(.a(new_n1389), .O(new_n1391));
  nor2 g01198(.a(new_n1391), .b(new_n1319), .O(new_n1392));
  nor2 g01199(.a(new_n1392), .b(new_n1390), .O(new_n1393));
  nor2 g01200(.a(new_n847), .b(new_n229), .O(new_n1394));
  inv1 g01201(.a(new_n1394), .O(new_n1395));
  nor2 g01202(.a(new_n1199), .b(new_n196), .O(new_n1396));
  nor2 g01203(.a(new_n1086), .b(new_n203), .O(new_n1397));
  nor2 g01204(.a(new_n1397), .b(new_n1396), .O(new_n1398));
  nor2 g01205(.a(new_n1199), .b(new_n203), .O(new_n1399));
  inv1 g01206(.a(new_n1399), .O(new_n1400));
  nor2 g01207(.a(new_n1400), .b(new_n1242), .O(new_n1401));
  nor2 g01208(.a(new_n1401), .b(new_n1398), .O(new_n1402));
  nor2 g01209(.a(new_n1402), .b(new_n1395), .O(new_n1403));
  inv1 g01210(.a(new_n1402), .O(new_n1404));
  nor2 g01211(.a(new_n1404), .b(new_n1394), .O(new_n1405));
  nor2 g01212(.a(new_n1405), .b(new_n1403), .O(new_n1406));
  nor2 g01213(.a(new_n1406), .b(new_n1393), .O(new_n1407));
  inv1 g01214(.a(new_n1393), .O(new_n1408));
  inv1 g01215(.a(new_n1406), .O(new_n1409));
  nor2 g01216(.a(new_n1409), .b(new_n1408), .O(new_n1410));
  nor2 g01217(.a(new_n1410), .b(new_n1407), .O(new_n1411));
  nor2 g01218(.a(new_n1411), .b(new_n1382), .O(new_n1412));
  inv1 g01219(.a(new_n1411), .O(new_n1413));
  nor2 g01220(.a(new_n1413), .b(new_n1381), .O(new_n1414));
  nor2 g01221(.a(new_n1414), .b(new_n1412), .O(new_n1415));
  nor2 g01222(.a(new_n1415), .b(new_n1370), .O(new_n1416));
  inv1 g01223(.a(new_n1370), .O(new_n1417));
  inv1 g01224(.a(new_n1415), .O(new_n1418));
  nor2 g01225(.a(new_n1418), .b(new_n1417), .O(new_n1419));
  nor2 g01226(.a(new_n1419), .b(new_n1416), .O(new_n1420));
  inv1 g01227(.a(new_n1420), .O(new_n1421));
  nor2 g01228(.a(new_n1288), .b(new_n1282), .O(new_n1422));
  inv1 g01229(.a(new_n1422), .O(new_n1423));
  inv1 g01230(.a(new_n1277), .O(new_n1424));
  inv1 g01231(.a(\a[21] ), .O(new_n1425));
  nor2 g01232(.a(new_n1425), .b(new_n198), .O(new_n1426));
  inv1 g01233(.a(new_n1426), .O(new_n1427));
  nor2 g01234(.a(new_n1427), .b(new_n1424), .O(new_n1428));
  nor2 g01235(.a(new_n1426), .b(new_n1277), .O(new_n1429));
  nor2 g01236(.a(new_n1429), .b(new_n1428), .O(new_n1430));
  inv1 g01237(.a(new_n1430), .O(new_n1431));
  nor2 g01238(.a(new_n1297), .b(new_n194), .O(new_n1432));
  inv1 g01239(.a(new_n1432), .O(new_n1433));
  nor2 g01240(.a(new_n1433), .b(new_n502), .O(new_n1434));
  nor2 g01241(.a(new_n1432), .b(\a[11] ), .O(new_n1435));
  nor2 g01242(.a(new_n1435), .b(new_n1434), .O(new_n1436));
  inv1 g01243(.a(new_n1436), .O(new_n1437));
  nor2 g01244(.a(new_n1437), .b(new_n1431), .O(new_n1438));
  nor2 g01245(.a(new_n1436), .b(new_n1430), .O(new_n1439));
  nor2 g01246(.a(new_n1439), .b(new_n1438), .O(new_n1440));
  nor2 g01247(.a(new_n1440), .b(new_n1423), .O(new_n1441));
  inv1 g01248(.a(new_n1440), .O(new_n1442));
  nor2 g01249(.a(new_n1442), .b(new_n1422), .O(new_n1443));
  nor2 g01250(.a(new_n1443), .b(new_n1441), .O(new_n1444));
  nor2 g01251(.a(new_n1327), .b(new_n1310), .O(new_n1445));
  inv1 g01252(.a(new_n1445), .O(new_n1446));
  nor2 g01253(.a(new_n1446), .b(new_n1444), .O(new_n1447));
  inv1 g01254(.a(new_n1444), .O(new_n1448));
  nor2 g01255(.a(new_n1445), .b(new_n1448), .O(new_n1449));
  nor2 g01256(.a(new_n1449), .b(new_n1447), .O(new_n1450));
  inv1 g01257(.a(new_n1450), .O(new_n1451));
  nor2 g01258(.a(new_n1332), .b(new_n1293), .O(new_n1452));
  nor2 g01259(.a(new_n1452), .b(new_n1451), .O(new_n1453));
  inv1 g01260(.a(new_n1452), .O(new_n1454));
  nor2 g01261(.a(new_n1454), .b(new_n1450), .O(new_n1455));
  nor2 g01262(.a(new_n1455), .b(new_n1453), .O(new_n1456));
  inv1 g01263(.a(new_n1456), .O(new_n1457));
  nor2 g01264(.a(new_n1457), .b(new_n1421), .O(new_n1458));
  nor2 g01265(.a(new_n1456), .b(new_n1420), .O(new_n1459));
  nor2 g01266(.a(new_n1459), .b(new_n1458), .O(new_n1460));
  inv1 g01267(.a(new_n1460), .O(new_n1461));
  nor2 g01268(.a(new_n1461), .b(new_n1351), .O(new_n1462));
  inv1 g01269(.a(new_n1351), .O(new_n1463));
  nor2 g01270(.a(new_n1460), .b(new_n1463), .O(new_n1464));
  nor2 g01271(.a(new_n1464), .b(new_n1462), .O(new_n1465));
  inv1 g01272(.a(new_n1465), .O(new_n1466));
  nor2 g01273(.a(new_n1346), .b(new_n1342), .O(new_n1467));
  nor2 g01274(.a(new_n1467), .b(new_n1466), .O(new_n1468));
  inv1 g01275(.a(new_n1467), .O(new_n1469));
  nor2 g01276(.a(new_n1469), .b(new_n1465), .O(new_n1470));
  nor2 g01277(.a(new_n1470), .b(new_n1468), .O(new_n1471));
  inv1 g01278(.a(new_n1471), .O(\asquared[22] ));
  nor2 g01279(.a(new_n1458), .b(new_n1453), .O(new_n1473));
  nor2 g01280(.a(new_n1405), .b(new_n1398), .O(new_n1474));
  nor2 g01281(.a(new_n1392), .b(new_n1385), .O(new_n1475));
  nor2 g01282(.a(new_n1475), .b(new_n1474), .O(new_n1476));
  inv1 g01283(.a(new_n1474), .O(new_n1477));
  inv1 g01284(.a(new_n1475), .O(new_n1478));
  nor2 g01285(.a(new_n1478), .b(new_n1477), .O(new_n1479));
  nor2 g01286(.a(new_n1479), .b(new_n1476), .O(new_n1480));
  nor2 g01287(.a(new_n1438), .b(new_n1428), .O(new_n1481));
  inv1 g01288(.a(new_n1481), .O(new_n1482));
  nor2 g01289(.a(new_n1482), .b(new_n1480), .O(new_n1483));
  inv1 g01290(.a(new_n1480), .O(new_n1484));
  nor2 g01291(.a(new_n1481), .b(new_n1484), .O(new_n1485));
  nor2 g01292(.a(new_n1485), .b(new_n1483), .O(new_n1486));
  nor2 g01293(.a(new_n1449), .b(new_n1443), .O(new_n1487));
  inv1 g01294(.a(new_n1487), .O(new_n1488));
  nor2 g01295(.a(new_n1488), .b(new_n1486), .O(new_n1489));
  inv1 g01296(.a(new_n1486), .O(new_n1490));
  nor2 g01297(.a(new_n1487), .b(new_n1490), .O(new_n1491));
  nor2 g01298(.a(new_n1491), .b(new_n1489), .O(new_n1492));
  inv1 g01299(.a(\a[22] ), .O(new_n1493));
  nor2 g01300(.a(new_n1493), .b(new_n198), .O(new_n1494));
  nor2 g01301(.a(new_n800), .b(new_n295), .O(new_n1495));
  nor2 g01302(.a(new_n1495), .b(new_n1386), .O(new_n1496));
  inv1 g01303(.a(new_n1384), .O(new_n1497));
  nor2 g01304(.a(new_n800), .b(new_n322), .O(new_n1498));
  inv1 g01305(.a(new_n1498), .O(new_n1499));
  nor2 g01306(.a(new_n1499), .b(new_n1497), .O(new_n1500));
  nor2 g01307(.a(new_n1500), .b(new_n1496), .O(new_n1501));
  inv1 g01308(.a(new_n1501), .O(new_n1502));
  nor2 g01309(.a(new_n1502), .b(new_n1494), .O(new_n1503));
  inv1 g01310(.a(new_n1494), .O(new_n1504));
  nor2 g01311(.a(new_n1501), .b(new_n1504), .O(new_n1505));
  nor2 g01312(.a(new_n1505), .b(new_n1503), .O(new_n1506));
  nor2 g01313(.a(new_n613), .b(new_n363), .O(new_n1507));
  inv1 g01314(.a(new_n1507), .O(new_n1508));
  nor2 g01315(.a(new_n1297), .b(new_n196), .O(new_n1509));
  nor2 g01316(.a(new_n1509), .b(new_n850), .O(new_n1510));
  inv1 g01317(.a(new_n1509), .O(new_n1511));
  nor2 g01318(.a(new_n1511), .b(new_n851), .O(new_n1512));
  nor2 g01319(.a(new_n1512), .b(new_n1510), .O(new_n1513));
  nor2 g01320(.a(new_n1513), .b(new_n1508), .O(new_n1514));
  inv1 g01321(.a(new_n1513), .O(new_n1515));
  nor2 g01322(.a(new_n1515), .b(new_n1507), .O(new_n1516));
  nor2 g01323(.a(new_n1516), .b(new_n1514), .O(new_n1517));
  nor2 g01324(.a(new_n1517), .b(new_n1506), .O(new_n1518));
  inv1 g01325(.a(new_n1506), .O(new_n1519));
  inv1 g01326(.a(new_n1517), .O(new_n1520));
  nor2 g01327(.a(new_n1520), .b(new_n1519), .O(new_n1521));
  nor2 g01328(.a(new_n1521), .b(new_n1518), .O(new_n1522));
  inv1 g01329(.a(new_n1522), .O(new_n1523));
  nor2 g01330(.a(new_n941), .b(new_n229), .O(new_n1524));
  nor2 g01331(.a(new_n1086), .b(new_n214), .O(new_n1525));
  nor2 g01332(.a(new_n1525), .b(new_n1524), .O(new_n1526));
  nor2 g01333(.a(new_n1086), .b(new_n229), .O(new_n1527));
  inv1 g01334(.a(new_n1527), .O(new_n1528));
  nor2 g01335(.a(new_n1528), .b(new_n1196), .O(new_n1529));
  nor2 g01336(.a(new_n1529), .b(new_n1526), .O(new_n1530));
  nor2 g01337(.a(new_n1530), .b(new_n1400), .O(new_n1531));
  inv1 g01338(.a(new_n1530), .O(new_n1532));
  nor2 g01339(.a(new_n1532), .b(new_n1399), .O(new_n1533));
  nor2 g01340(.a(new_n1533), .b(new_n1531), .O(new_n1534));
  nor2 g01341(.a(new_n1534), .b(new_n1523), .O(new_n1535));
  inv1 g01342(.a(new_n1534), .O(new_n1536));
  nor2 g01343(.a(new_n1536), .b(new_n1522), .O(new_n1537));
  nor2 g01344(.a(new_n1537), .b(new_n1535), .O(new_n1538));
  nor2 g01345(.a(new_n1538), .b(new_n1492), .O(new_n1539));
  inv1 g01346(.a(new_n1492), .O(new_n1540));
  inv1 g01347(.a(new_n1538), .O(new_n1541));
  nor2 g01348(.a(new_n1541), .b(new_n1540), .O(new_n1542));
  nor2 g01349(.a(new_n1542), .b(new_n1539), .O(new_n1543));
  inv1 g01350(.a(new_n1543), .O(new_n1544));
  nor2 g01351(.a(new_n1419), .b(new_n1369), .O(new_n1545));
  nor2 g01352(.a(new_n1363), .b(new_n1357), .O(new_n1546));
  inv1 g01353(.a(new_n1434), .O(new_n1547));
  nor2 g01354(.a(new_n1425), .b(new_n194), .O(new_n1548));
  nor2 g01355(.a(new_n1548), .b(new_n1374), .O(new_n1549));
  inv1 g01356(.a(new_n1548), .O(new_n1550));
  nor2 g01357(.a(new_n1550), .b(new_n1375), .O(new_n1551));
  nor2 g01358(.a(new_n1551), .b(new_n1549), .O(new_n1552));
  inv1 g01359(.a(new_n1552), .O(new_n1553));
  nor2 g01360(.a(new_n1553), .b(new_n1547), .O(new_n1554));
  nor2 g01361(.a(new_n1552), .b(new_n1434), .O(new_n1555));
  nor2 g01362(.a(new_n1555), .b(new_n1554), .O(new_n1556));
  inv1 g01363(.a(new_n1556), .O(new_n1557));
  nor2 g01364(.a(new_n1380), .b(new_n1373), .O(new_n1558));
  inv1 g01365(.a(new_n1558), .O(new_n1559));
  nor2 g01366(.a(new_n1559), .b(new_n1557), .O(new_n1560));
  nor2 g01367(.a(new_n1558), .b(new_n1556), .O(new_n1561));
  nor2 g01368(.a(new_n1561), .b(new_n1560), .O(new_n1562));
  inv1 g01369(.a(new_n1562), .O(new_n1563));
  nor2 g01370(.a(new_n1563), .b(new_n1546), .O(new_n1564));
  inv1 g01371(.a(new_n1546), .O(new_n1565));
  nor2 g01372(.a(new_n1562), .b(new_n1565), .O(new_n1566));
  nor2 g01373(.a(new_n1566), .b(new_n1564), .O(new_n1567));
  inv1 g01374(.a(new_n1567), .O(new_n1568));
  nor2 g01375(.a(new_n1414), .b(new_n1407), .O(new_n1569));
  nor2 g01376(.a(new_n1569), .b(new_n1568), .O(new_n1570));
  inv1 g01377(.a(new_n1569), .O(new_n1571));
  nor2 g01378(.a(new_n1571), .b(new_n1567), .O(new_n1572));
  nor2 g01379(.a(new_n1572), .b(new_n1570), .O(new_n1573));
  inv1 g01380(.a(new_n1573), .O(new_n1574));
  nor2 g01381(.a(new_n1574), .b(new_n1545), .O(new_n1575));
  inv1 g01382(.a(new_n1545), .O(new_n1576));
  nor2 g01383(.a(new_n1573), .b(new_n1576), .O(new_n1577));
  nor2 g01384(.a(new_n1577), .b(new_n1575), .O(new_n1578));
  inv1 g01385(.a(new_n1578), .O(new_n1579));
  nor2 g01386(.a(new_n1579), .b(new_n1544), .O(new_n1580));
  nor2 g01387(.a(new_n1578), .b(new_n1543), .O(new_n1581));
  nor2 g01388(.a(new_n1581), .b(new_n1580), .O(new_n1582));
  inv1 g01389(.a(new_n1582), .O(new_n1583));
  nor2 g01390(.a(new_n1583), .b(new_n1473), .O(new_n1584));
  inv1 g01391(.a(new_n1473), .O(new_n1585));
  nor2 g01392(.a(new_n1582), .b(new_n1585), .O(new_n1586));
  nor2 g01393(.a(new_n1586), .b(new_n1584), .O(new_n1587));
  inv1 g01394(.a(new_n1587), .O(new_n1588));
  nor2 g01395(.a(new_n1468), .b(new_n1464), .O(new_n1589));
  nor2 g01396(.a(new_n1589), .b(new_n1588), .O(new_n1590));
  inv1 g01397(.a(new_n1589), .O(new_n1591));
  nor2 g01398(.a(new_n1591), .b(new_n1587), .O(new_n1592));
  nor2 g01399(.a(new_n1592), .b(new_n1590), .O(new_n1593));
  inv1 g01400(.a(new_n1593), .O(\asquared[23] ));
  nor2 g01401(.a(new_n1580), .b(new_n1575), .O(new_n1595));
  inv1 g01402(.a(new_n1595), .O(new_n1596));
  nor2 g01403(.a(new_n1570), .b(new_n1564), .O(new_n1597));
  nor2 g01404(.a(new_n1560), .b(new_n1554), .O(new_n1598));
  inv1 g01405(.a(new_n1598), .O(new_n1599));
  nor2 g01406(.a(new_n941), .b(new_n257), .O(new_n1600));
  nor2 g01407(.a(new_n1297), .b(new_n203), .O(new_n1601));
  nor2 g01408(.a(new_n1601), .b(new_n1527), .O(new_n1602));
  inv1 g01409(.a(new_n1397), .O(new_n1603));
  nor2 g01410(.a(new_n1297), .b(new_n229), .O(new_n1604));
  inv1 g01411(.a(new_n1604), .O(new_n1605));
  nor2 g01412(.a(new_n1605), .b(new_n1603), .O(new_n1606));
  nor2 g01413(.a(new_n1606), .b(new_n1602), .O(new_n1607));
  inv1 g01414(.a(new_n1607), .O(new_n1608));
  nor2 g01415(.a(new_n1608), .b(new_n1600), .O(new_n1609));
  inv1 g01416(.a(new_n1600), .O(new_n1610));
  nor2 g01417(.a(new_n1607), .b(new_n1610), .O(new_n1611));
  nor2 g01418(.a(new_n1611), .b(new_n1609), .O(new_n1612));
  nor2 g01419(.a(new_n1199), .b(new_n214), .O(new_n1613));
  inv1 g01420(.a(new_n1613), .O(new_n1614));
  nor2 g01421(.a(new_n569), .b(new_n502), .O(new_n1615));
  nor2 g01422(.a(new_n613), .b(new_n438), .O(new_n1616));
  nor2 g01423(.a(new_n1616), .b(new_n1615), .O(new_n1617));
  nor2 g01424(.a(new_n613), .b(new_n502), .O(new_n1618));
  inv1 g01425(.a(new_n1618), .O(new_n1619));
  nor2 g01426(.a(new_n1619), .b(new_n1375), .O(new_n1620));
  nor2 g01427(.a(new_n1620), .b(new_n1617), .O(new_n1621));
  nor2 g01428(.a(new_n1621), .b(new_n1614), .O(new_n1622));
  inv1 g01429(.a(new_n1621), .O(new_n1623));
  nor2 g01430(.a(new_n1623), .b(new_n1613), .O(new_n1624));
  nor2 g01431(.a(new_n1624), .b(new_n1622), .O(new_n1625));
  nor2 g01432(.a(new_n1625), .b(new_n1612), .O(new_n1626));
  inv1 g01433(.a(new_n1612), .O(new_n1627));
  inv1 g01434(.a(new_n1625), .O(new_n1628));
  nor2 g01435(.a(new_n1628), .b(new_n1627), .O(new_n1629));
  nor2 g01436(.a(new_n1629), .b(new_n1626), .O(new_n1630));
  nor2 g01437(.a(new_n1630), .b(new_n1599), .O(new_n1631));
  inv1 g01438(.a(new_n1630), .O(new_n1632));
  nor2 g01439(.a(new_n1632), .b(new_n1598), .O(new_n1633));
  nor2 g01440(.a(new_n1633), .b(new_n1631), .O(new_n1634));
  nor2 g01441(.a(new_n847), .b(new_n295), .O(new_n1635));
  inv1 g01442(.a(new_n1635), .O(new_n1636));
  nor2 g01443(.a(new_n699), .b(new_n363), .O(new_n1637));
  nor2 g01444(.a(new_n1637), .b(new_n1498), .O(new_n1638));
  nor2 g01445(.a(new_n800), .b(new_n363), .O(new_n1639));
  inv1 g01446(.a(new_n1639), .O(new_n1640));
  nor2 g01447(.a(new_n1640), .b(new_n1387), .O(new_n1641));
  nor2 g01448(.a(new_n1641), .b(new_n1638), .O(new_n1642));
  nor2 g01449(.a(new_n1642), .b(new_n1636), .O(new_n1643));
  inv1 g01450(.a(new_n1642), .O(new_n1644));
  nor2 g01451(.a(new_n1644), .b(new_n1635), .O(new_n1645));
  nor2 g01452(.a(new_n1645), .b(new_n1643), .O(new_n1646));
  inv1 g01453(.a(\a[23] ), .O(new_n1647));
  nor2 g01454(.a(new_n1647), .b(new_n198), .O(new_n1648));
  nor2 g01455(.a(new_n1425), .b(new_n196), .O(new_n1649));
  nor2 g01456(.a(new_n1649), .b(new_n1648), .O(new_n1650));
  nor2 g01457(.a(new_n1647), .b(new_n196), .O(new_n1651));
  inv1 g01458(.a(new_n1651), .O(new_n1652));
  nor2 g01459(.a(new_n1652), .b(new_n1427), .O(new_n1653));
  nor2 g01460(.a(new_n1653), .b(new_n1650), .O(new_n1654));
  inv1 g01461(.a(new_n1654), .O(new_n1655));
  nor2 g01462(.a(new_n1655), .b(new_n1551), .O(new_n1656));
  inv1 g01463(.a(new_n1551), .O(new_n1657));
  nor2 g01464(.a(new_n1654), .b(new_n1657), .O(new_n1658));
  nor2 g01465(.a(new_n1658), .b(new_n1656), .O(new_n1659));
  nor2 g01466(.a(new_n1503), .b(new_n1496), .O(new_n1660));
  inv1 g01467(.a(new_n1660), .O(new_n1661));
  nor2 g01468(.a(new_n1661), .b(new_n1659), .O(new_n1662));
  inv1 g01469(.a(new_n1659), .O(new_n1663));
  nor2 g01470(.a(new_n1660), .b(new_n1663), .O(new_n1664));
  nor2 g01471(.a(new_n1664), .b(new_n1662), .O(new_n1665));
  inv1 g01472(.a(new_n1665), .O(new_n1666));
  nor2 g01473(.a(new_n1666), .b(new_n1646), .O(new_n1667));
  inv1 g01474(.a(new_n1646), .O(new_n1668));
  nor2 g01475(.a(new_n1665), .b(new_n1668), .O(new_n1669));
  nor2 g01476(.a(new_n1669), .b(new_n1667), .O(new_n1670));
  nor2 g01477(.a(new_n1670), .b(new_n1634), .O(new_n1671));
  inv1 g01478(.a(new_n1634), .O(new_n1672));
  inv1 g01479(.a(new_n1670), .O(new_n1673));
  nor2 g01480(.a(new_n1673), .b(new_n1672), .O(new_n1674));
  nor2 g01481(.a(new_n1674), .b(new_n1671), .O(new_n1675));
  inv1 g01482(.a(new_n1675), .O(new_n1676));
  nor2 g01483(.a(new_n1676), .b(new_n1597), .O(new_n1677));
  inv1 g01484(.a(new_n1597), .O(new_n1678));
  nor2 g01485(.a(new_n1675), .b(new_n1678), .O(new_n1679));
  nor2 g01486(.a(new_n1679), .b(new_n1677), .O(new_n1680));
  inv1 g01487(.a(new_n1680), .O(new_n1681));
  nor2 g01488(.a(new_n1542), .b(new_n1491), .O(new_n1682));
  nor2 g01489(.a(new_n1485), .b(new_n1479), .O(new_n1683));
  inv1 g01490(.a(new_n1683), .O(new_n1684));
  nor2 g01491(.a(new_n1535), .b(new_n1518), .O(new_n1685));
  inv1 g01492(.a(new_n1685), .O(new_n1686));
  nor2 g01493(.a(new_n1686), .b(new_n1684), .O(new_n1687));
  nor2 g01494(.a(new_n1685), .b(new_n1683), .O(new_n1688));
  nor2 g01495(.a(new_n1688), .b(new_n1687), .O(new_n1689));
  inv1 g01496(.a(new_n1689), .O(new_n1690));
  nor2 g01497(.a(new_n1493), .b(new_n194), .O(new_n1691));
  inv1 g01498(.a(new_n1691), .O(new_n1692));
  nor2 g01499(.a(new_n1692), .b(new_n569), .O(new_n1693));
  nor2 g01500(.a(new_n1691), .b(\a[12] ), .O(new_n1694));
  nor2 g01501(.a(new_n1694), .b(new_n1693), .O(new_n1695));
  nor2 g01502(.a(new_n1533), .b(new_n1526), .O(new_n1696));
  nor2 g01503(.a(new_n1696), .b(new_n1695), .O(new_n1697));
  inv1 g01504(.a(new_n1695), .O(new_n1698));
  inv1 g01505(.a(new_n1696), .O(new_n1699));
  nor2 g01506(.a(new_n1699), .b(new_n1698), .O(new_n1700));
  nor2 g01507(.a(new_n1700), .b(new_n1697), .O(new_n1701));
  inv1 g01508(.a(new_n1701), .O(new_n1702));
  nor2 g01509(.a(new_n1516), .b(new_n1510), .O(new_n1703));
  inv1 g01510(.a(new_n1703), .O(new_n1704));
  nor2 g01511(.a(new_n1704), .b(new_n1702), .O(new_n1705));
  nor2 g01512(.a(new_n1703), .b(new_n1701), .O(new_n1706));
  nor2 g01513(.a(new_n1706), .b(new_n1705), .O(new_n1707));
  inv1 g01514(.a(new_n1707), .O(new_n1708));
  nor2 g01515(.a(new_n1708), .b(new_n1690), .O(new_n1709));
  nor2 g01516(.a(new_n1707), .b(new_n1689), .O(new_n1710));
  nor2 g01517(.a(new_n1710), .b(new_n1709), .O(new_n1711));
  inv1 g01518(.a(new_n1711), .O(new_n1712));
  nor2 g01519(.a(new_n1712), .b(new_n1682), .O(new_n1713));
  inv1 g01520(.a(new_n1682), .O(new_n1714));
  nor2 g01521(.a(new_n1711), .b(new_n1714), .O(new_n1715));
  nor2 g01522(.a(new_n1715), .b(new_n1713), .O(new_n1716));
  inv1 g01523(.a(new_n1716), .O(new_n1717));
  nor2 g01524(.a(new_n1717), .b(new_n1681), .O(new_n1718));
  nor2 g01525(.a(new_n1716), .b(new_n1680), .O(new_n1719));
  nor2 g01526(.a(new_n1719), .b(new_n1718), .O(new_n1720));
  nor2 g01527(.a(new_n1720), .b(new_n1596), .O(new_n1721));
  inv1 g01528(.a(new_n1720), .O(new_n1722));
  nor2 g01529(.a(new_n1722), .b(new_n1595), .O(new_n1723));
  nor2 g01530(.a(new_n1723), .b(new_n1721), .O(new_n1724));
  inv1 g01531(.a(new_n1724), .O(new_n1725));
  nor2 g01532(.a(new_n1590), .b(new_n1586), .O(new_n1726));
  nor2 g01533(.a(new_n1726), .b(new_n1725), .O(new_n1727));
  inv1 g01534(.a(new_n1726), .O(new_n1728));
  nor2 g01535(.a(new_n1728), .b(new_n1724), .O(new_n1729));
  nor2 g01536(.a(new_n1729), .b(new_n1727), .O(new_n1730));
  inv1 g01537(.a(new_n1730), .O(\asquared[24] ));
  nor2 g01538(.a(new_n1718), .b(new_n1713), .O(new_n1732));
  nor2 g01539(.a(new_n1705), .b(new_n1700), .O(new_n1733));
  inv1 g01540(.a(new_n1733), .O(new_n1734));
  inv1 g01541(.a(new_n1693), .O(new_n1735));
  inv1 g01542(.a(\a[24] ), .O(new_n1736));
  nor2 g01543(.a(new_n1736), .b(new_n198), .O(new_n1737));
  inv1 g01544(.a(new_n1737), .O(new_n1738));
  nor2 g01545(.a(new_n1738), .b(new_n1735), .O(new_n1739));
  nor2 g01546(.a(new_n1737), .b(new_n1693), .O(new_n1740));
  nor2 g01547(.a(new_n1740), .b(new_n1739), .O(new_n1741));
  inv1 g01548(.a(new_n1741), .O(new_n1742));
  nor2 g01549(.a(new_n1647), .b(new_n194), .O(new_n1743));
  nor2 g01550(.a(new_n1743), .b(new_n1618), .O(new_n1744));
  inv1 g01551(.a(new_n1743), .O(new_n1745));
  nor2 g01552(.a(new_n1745), .b(new_n1619), .O(new_n1746));
  nor2 g01553(.a(new_n1746), .b(new_n1744), .O(new_n1747));
  inv1 g01554(.a(new_n1747), .O(new_n1748));
  nor2 g01555(.a(new_n1748), .b(new_n1742), .O(new_n1749));
  nor2 g01556(.a(new_n1747), .b(new_n1741), .O(new_n1750));
  nor2 g01557(.a(new_n1750), .b(new_n1749), .O(new_n1751));
  inv1 g01558(.a(new_n1751), .O(new_n1752));
  nor2 g01559(.a(new_n941), .b(new_n295), .O(new_n1753));
  inv1 g01560(.a(new_n1753), .O(new_n1754));
  nor2 g01561(.a(new_n1493), .b(new_n196), .O(new_n1755));
  nor2 g01562(.a(new_n1086), .b(new_n257), .O(new_n1756));
  nor2 g01563(.a(new_n1756), .b(new_n1755), .O(new_n1757));
  nor2 g01564(.a(new_n1493), .b(new_n257), .O(new_n1758));
  inv1 g01565(.a(new_n1758), .O(new_n1759));
  nor2 g01566(.a(new_n1759), .b(new_n1242), .O(new_n1760));
  nor2 g01567(.a(new_n1760), .b(new_n1757), .O(new_n1761));
  nor2 g01568(.a(new_n1761), .b(new_n1754), .O(new_n1762));
  inv1 g01569(.a(new_n1761), .O(new_n1763));
  nor2 g01570(.a(new_n1763), .b(new_n1753), .O(new_n1764));
  nor2 g01571(.a(new_n1764), .b(new_n1762), .O(new_n1765));
  nor2 g01572(.a(new_n1765), .b(new_n1752), .O(new_n1766));
  inv1 g01573(.a(new_n1765), .O(new_n1767));
  nor2 g01574(.a(new_n1767), .b(new_n1751), .O(new_n1768));
  nor2 g01575(.a(new_n1768), .b(new_n1766), .O(new_n1769));
  nor2 g01576(.a(new_n1769), .b(new_n1734), .O(new_n1770));
  inv1 g01577(.a(new_n1769), .O(new_n1771));
  nor2 g01578(.a(new_n1771), .b(new_n1733), .O(new_n1772));
  nor2 g01579(.a(new_n1772), .b(new_n1770), .O(new_n1773));
  nor2 g01580(.a(new_n847), .b(new_n322), .O(new_n1774));
  inv1 g01581(.a(new_n1774), .O(new_n1775));
  nor2 g01582(.a(new_n699), .b(new_n438), .O(new_n1776));
  nor2 g01583(.a(new_n1776), .b(new_n1639), .O(new_n1777));
  inv1 g01584(.a(new_n1637), .O(new_n1778));
  nor2 g01585(.a(new_n800), .b(new_n438), .O(new_n1779));
  inv1 g01586(.a(new_n1779), .O(new_n1780));
  nor2 g01587(.a(new_n1780), .b(new_n1778), .O(new_n1781));
  nor2 g01588(.a(new_n1781), .b(new_n1777), .O(new_n1782));
  nor2 g01589(.a(new_n1782), .b(new_n1775), .O(new_n1783));
  inv1 g01590(.a(new_n1782), .O(new_n1784));
  nor2 g01591(.a(new_n1784), .b(new_n1774), .O(new_n1785));
  nor2 g01592(.a(new_n1785), .b(new_n1783), .O(new_n1786));
  nor2 g01593(.a(new_n1425), .b(new_n203), .O(new_n1787));
  inv1 g01594(.a(new_n1787), .O(new_n1788));
  nor2 g01595(.a(new_n1199), .b(new_n229), .O(new_n1789));
  nor2 g01596(.a(new_n1297), .b(new_n214), .O(new_n1790));
  nor2 g01597(.a(new_n1790), .b(new_n1789), .O(new_n1791));
  nor2 g01598(.a(new_n1614), .b(new_n1605), .O(new_n1792));
  nor2 g01599(.a(new_n1792), .b(new_n1791), .O(new_n1793));
  nor2 g01600(.a(new_n1793), .b(new_n1788), .O(new_n1794));
  inv1 g01601(.a(new_n1793), .O(new_n1795));
  nor2 g01602(.a(new_n1795), .b(new_n1787), .O(new_n1796));
  nor2 g01603(.a(new_n1796), .b(new_n1794), .O(new_n1797));
  nor2 g01604(.a(new_n1656), .b(new_n1650), .O(new_n1798));
  inv1 g01605(.a(new_n1798), .O(new_n1799));
  nor2 g01606(.a(new_n1799), .b(new_n1797), .O(new_n1800));
  inv1 g01607(.a(new_n1797), .O(new_n1801));
  nor2 g01608(.a(new_n1798), .b(new_n1801), .O(new_n1802));
  nor2 g01609(.a(new_n1802), .b(new_n1800), .O(new_n1803));
  inv1 g01610(.a(new_n1803), .O(new_n1804));
  nor2 g01611(.a(new_n1804), .b(new_n1786), .O(new_n1805));
  inv1 g01612(.a(new_n1786), .O(new_n1806));
  nor2 g01613(.a(new_n1803), .b(new_n1806), .O(new_n1807));
  nor2 g01614(.a(new_n1807), .b(new_n1805), .O(new_n1808));
  nor2 g01615(.a(new_n1808), .b(new_n1773), .O(new_n1809));
  inv1 g01616(.a(new_n1773), .O(new_n1810));
  inv1 g01617(.a(new_n1808), .O(new_n1811));
  nor2 g01618(.a(new_n1811), .b(new_n1810), .O(new_n1812));
  nor2 g01619(.a(new_n1812), .b(new_n1809), .O(new_n1813));
  inv1 g01620(.a(new_n1813), .O(new_n1814));
  nor2 g01621(.a(new_n1709), .b(new_n1688), .O(new_n1815));
  nor2 g01622(.a(new_n1815), .b(new_n1814), .O(new_n1816));
  inv1 g01623(.a(new_n1815), .O(new_n1817));
  nor2 g01624(.a(new_n1817), .b(new_n1813), .O(new_n1818));
  nor2 g01625(.a(new_n1818), .b(new_n1816), .O(new_n1819));
  inv1 g01626(.a(new_n1819), .O(new_n1820));
  nor2 g01627(.a(new_n1677), .b(new_n1674), .O(new_n1821));
  nor2 g01628(.a(new_n1624), .b(new_n1617), .O(new_n1822));
  nor2 g01629(.a(new_n1609), .b(new_n1602), .O(new_n1823));
  nor2 g01630(.a(new_n1823), .b(new_n1822), .O(new_n1824));
  inv1 g01631(.a(new_n1822), .O(new_n1825));
  inv1 g01632(.a(new_n1823), .O(new_n1826));
  nor2 g01633(.a(new_n1826), .b(new_n1825), .O(new_n1827));
  nor2 g01634(.a(new_n1827), .b(new_n1824), .O(new_n1828));
  nor2 g01635(.a(new_n1645), .b(new_n1638), .O(new_n1829));
  nor2 g01636(.a(new_n1829), .b(new_n1828), .O(new_n1830));
  inv1 g01637(.a(new_n1828), .O(new_n1831));
  inv1 g01638(.a(new_n1829), .O(new_n1832));
  nor2 g01639(.a(new_n1832), .b(new_n1831), .O(new_n1833));
  nor2 g01640(.a(new_n1833), .b(new_n1830), .O(new_n1834));
  inv1 g01641(.a(new_n1834), .O(new_n1835));
  nor2 g01642(.a(new_n1633), .b(new_n1626), .O(new_n1836));
  inv1 g01643(.a(new_n1836), .O(new_n1837));
  nor2 g01644(.a(new_n1667), .b(new_n1662), .O(new_n1838));
  inv1 g01645(.a(new_n1838), .O(new_n1839));
  nor2 g01646(.a(new_n1839), .b(new_n1837), .O(new_n1840));
  nor2 g01647(.a(new_n1838), .b(new_n1836), .O(new_n1841));
  nor2 g01648(.a(new_n1841), .b(new_n1840), .O(new_n1842));
  inv1 g01649(.a(new_n1842), .O(new_n1843));
  nor2 g01650(.a(new_n1843), .b(new_n1835), .O(new_n1844));
  nor2 g01651(.a(new_n1842), .b(new_n1834), .O(new_n1845));
  nor2 g01652(.a(new_n1845), .b(new_n1844), .O(new_n1846));
  inv1 g01653(.a(new_n1846), .O(new_n1847));
  nor2 g01654(.a(new_n1847), .b(new_n1821), .O(new_n1848));
  inv1 g01655(.a(new_n1821), .O(new_n1849));
  nor2 g01656(.a(new_n1846), .b(new_n1849), .O(new_n1850));
  nor2 g01657(.a(new_n1850), .b(new_n1848), .O(new_n1851));
  inv1 g01658(.a(new_n1851), .O(new_n1852));
  nor2 g01659(.a(new_n1852), .b(new_n1820), .O(new_n1853));
  nor2 g01660(.a(new_n1851), .b(new_n1819), .O(new_n1854));
  nor2 g01661(.a(new_n1854), .b(new_n1853), .O(new_n1855));
  inv1 g01662(.a(new_n1855), .O(new_n1856));
  nor2 g01663(.a(new_n1856), .b(new_n1732), .O(new_n1857));
  inv1 g01664(.a(new_n1732), .O(new_n1858));
  nor2 g01665(.a(new_n1855), .b(new_n1858), .O(new_n1859));
  nor2 g01666(.a(new_n1859), .b(new_n1857), .O(new_n1860));
  inv1 g01667(.a(new_n1860), .O(new_n1861));
  nor2 g01668(.a(new_n1727), .b(new_n1721), .O(new_n1862));
  nor2 g01669(.a(new_n1862), .b(new_n1861), .O(new_n1863));
  inv1 g01670(.a(new_n1862), .O(new_n1864));
  nor2 g01671(.a(new_n1864), .b(new_n1860), .O(new_n1865));
  nor2 g01672(.a(new_n1865), .b(new_n1863), .O(new_n1866));
  inv1 g01673(.a(new_n1866), .O(\asquared[25] ));
  nor2 g01674(.a(new_n1853), .b(new_n1848), .O(new_n1868));
  inv1 g01675(.a(new_n1868), .O(new_n1869));
  nor2 g01676(.a(new_n1764), .b(new_n1757), .O(new_n1870));
  nor2 g01677(.a(new_n1785), .b(new_n1777), .O(new_n1871));
  nor2 g01678(.a(new_n1871), .b(new_n1870), .O(new_n1872));
  inv1 g01679(.a(new_n1870), .O(new_n1873));
  inv1 g01680(.a(new_n1871), .O(new_n1874));
  nor2 g01681(.a(new_n1874), .b(new_n1873), .O(new_n1875));
  nor2 g01682(.a(new_n1875), .b(new_n1872), .O(new_n1876));
  nor2 g01683(.a(new_n1749), .b(new_n1739), .O(new_n1877));
  inv1 g01684(.a(new_n1877), .O(new_n1878));
  nor2 g01685(.a(new_n1878), .b(new_n1876), .O(new_n1879));
  inv1 g01686(.a(new_n1876), .O(new_n1880));
  nor2 g01687(.a(new_n1877), .b(new_n1880), .O(new_n1881));
  nor2 g01688(.a(new_n1881), .b(new_n1879), .O(new_n1882));
  nor2 g01689(.a(new_n1805), .b(new_n1800), .O(new_n1883));
  inv1 g01690(.a(new_n1883), .O(new_n1884));
  nor2 g01691(.a(new_n1884), .b(new_n1882), .O(new_n1885));
  inv1 g01692(.a(new_n1882), .O(new_n1886));
  nor2 g01693(.a(new_n1883), .b(new_n1886), .O(new_n1887));
  nor2 g01694(.a(new_n1887), .b(new_n1885), .O(new_n1888));
  nor2 g01695(.a(new_n1772), .b(new_n1766), .O(new_n1889));
  inv1 g01696(.a(new_n1889), .O(new_n1890));
  nor2 g01697(.a(new_n1890), .b(new_n1888), .O(new_n1891));
  inv1 g01698(.a(new_n1888), .O(new_n1892));
  nor2 g01699(.a(new_n1889), .b(new_n1892), .O(new_n1893));
  nor2 g01700(.a(new_n1893), .b(new_n1891), .O(new_n1894));
  inv1 g01701(.a(new_n1894), .O(new_n1895));
  nor2 g01702(.a(new_n1816), .b(new_n1812), .O(new_n1896));
  nor2 g01703(.a(new_n1896), .b(new_n1895), .O(new_n1897));
  inv1 g01704(.a(new_n1896), .O(new_n1898));
  nor2 g01705(.a(new_n1898), .b(new_n1894), .O(new_n1899));
  nor2 g01706(.a(new_n1899), .b(new_n1897), .O(new_n1900));
  inv1 g01707(.a(new_n1900), .O(new_n1901));
  nor2 g01708(.a(new_n1844), .b(new_n1841), .O(new_n1902));
  inv1 g01709(.a(\a[25] ), .O(new_n1903));
  nor2 g01710(.a(new_n1903), .b(new_n198), .O(new_n1904));
  nor2 g01711(.a(new_n1904), .b(new_n1651), .O(new_n1905));
  inv1 g01712(.a(new_n1648), .O(new_n1906));
  nor2 g01713(.a(new_n1903), .b(new_n196), .O(new_n1907));
  inv1 g01714(.a(new_n1907), .O(new_n1908));
  nor2 g01715(.a(new_n1908), .b(new_n1906), .O(new_n1909));
  nor2 g01716(.a(new_n1909), .b(new_n1905), .O(new_n1910));
  inv1 g01717(.a(new_n1910), .O(new_n1911));
  nor2 g01718(.a(new_n1911), .b(new_n1779), .O(new_n1912));
  nor2 g01719(.a(new_n1910), .b(new_n1780), .O(new_n1913));
  nor2 g01720(.a(new_n1913), .b(new_n1912), .O(new_n1914));
  nor2 g01721(.a(new_n1086), .b(new_n295), .O(new_n1915));
  inv1 g01722(.a(new_n1915), .O(new_n1916));
  nor2 g01723(.a(new_n941), .b(new_n322), .O(new_n1917));
  nor2 g01724(.a(new_n1917), .b(new_n988), .O(new_n1918));
  nor2 g01725(.a(new_n941), .b(new_n363), .O(new_n1919));
  inv1 g01726(.a(new_n1919), .O(new_n1920));
  nor2 g01727(.a(new_n1920), .b(new_n1775), .O(new_n1921));
  nor2 g01728(.a(new_n1921), .b(new_n1918), .O(new_n1922));
  nor2 g01729(.a(new_n1922), .b(new_n1916), .O(new_n1923));
  inv1 g01730(.a(new_n1922), .O(new_n1924));
  nor2 g01731(.a(new_n1924), .b(new_n1915), .O(new_n1925));
  nor2 g01732(.a(new_n1925), .b(new_n1923), .O(new_n1926));
  nor2 g01733(.a(new_n1926), .b(new_n1914), .O(new_n1927));
  inv1 g01734(.a(new_n1914), .O(new_n1928));
  inv1 g01735(.a(new_n1926), .O(new_n1929));
  nor2 g01736(.a(new_n1929), .b(new_n1928), .O(new_n1930));
  nor2 g01737(.a(new_n1930), .b(new_n1927), .O(new_n1931));
  nor2 g01738(.a(new_n1199), .b(new_n257), .O(new_n1932));
  inv1 g01739(.a(new_n1932), .O(new_n1933));
  nor2 g01740(.a(new_n1493), .b(new_n203), .O(new_n1934));
  nor2 g01741(.a(new_n1425), .b(new_n214), .O(new_n1935));
  nor2 g01742(.a(new_n1935), .b(new_n1934), .O(new_n1936));
  nor2 g01743(.a(new_n1493), .b(new_n214), .O(new_n1937));
  inv1 g01744(.a(new_n1937), .O(new_n1938));
  nor2 g01745(.a(new_n1938), .b(new_n1788), .O(new_n1939));
  nor2 g01746(.a(new_n1939), .b(new_n1936), .O(new_n1940));
  nor2 g01747(.a(new_n1940), .b(new_n1933), .O(new_n1941));
  inv1 g01748(.a(new_n1940), .O(new_n1942));
  nor2 g01749(.a(new_n1942), .b(new_n1932), .O(new_n1943));
  nor2 g01750(.a(new_n1943), .b(new_n1941), .O(new_n1944));
  inv1 g01751(.a(new_n1944), .O(new_n1945));
  nor2 g01752(.a(new_n1945), .b(new_n1931), .O(new_n1946));
  inv1 g01753(.a(new_n1931), .O(new_n1947));
  nor2 g01754(.a(new_n1944), .b(new_n1947), .O(new_n1948));
  nor2 g01755(.a(new_n1948), .b(new_n1946), .O(new_n1949));
  inv1 g01756(.a(new_n1949), .O(new_n1950));
  nor2 g01757(.a(new_n1950), .b(new_n1902), .O(new_n1951));
  inv1 g01758(.a(new_n1902), .O(new_n1952));
  nor2 g01759(.a(new_n1949), .b(new_n1952), .O(new_n1953));
  nor2 g01760(.a(new_n1953), .b(new_n1951), .O(new_n1954));
  inv1 g01761(.a(new_n1954), .O(new_n1955));
  nor2 g01762(.a(new_n1736), .b(new_n194), .O(new_n1956));
  inv1 g01763(.a(new_n1956), .O(new_n1957));
  nor2 g01764(.a(new_n1746), .b(new_n613), .O(new_n1958));
  nor2 g01765(.a(new_n1958), .b(new_n1957), .O(new_n1959));
  inv1 g01766(.a(new_n1958), .O(new_n1960));
  nor2 g01767(.a(new_n1960), .b(new_n1956), .O(new_n1961));
  nor2 g01768(.a(new_n1961), .b(new_n1959), .O(new_n1962));
  nor2 g01769(.a(new_n1796), .b(new_n1791), .O(new_n1963));
  inv1 g01770(.a(new_n1963), .O(new_n1964));
  nor2 g01771(.a(new_n1964), .b(new_n1962), .O(new_n1965));
  inv1 g01772(.a(new_n1962), .O(new_n1966));
  nor2 g01773(.a(new_n1963), .b(new_n1966), .O(new_n1967));
  nor2 g01774(.a(new_n1967), .b(new_n1965), .O(new_n1968));
  inv1 g01775(.a(new_n1968), .O(new_n1969));
  nor2 g01776(.a(new_n1833), .b(new_n1827), .O(new_n1970));
  nor2 g01777(.a(new_n613), .b(new_n569), .O(new_n1971));
  nor2 g01778(.a(new_n699), .b(new_n502), .O(new_n1972));
  nor2 g01779(.a(new_n1972), .b(new_n1971), .O(new_n1973));
  inv1 g01780(.a(new_n1971), .O(new_n1974));
  inv1 g01781(.a(new_n1972), .O(new_n1975));
  nor2 g01782(.a(new_n1975), .b(new_n1974), .O(new_n1976));
  nor2 g01783(.a(new_n1976), .b(new_n1973), .O(new_n1977));
  nor2 g01784(.a(new_n1977), .b(new_n1605), .O(new_n1978));
  inv1 g01785(.a(new_n1977), .O(new_n1979));
  nor2 g01786(.a(new_n1979), .b(new_n1604), .O(new_n1980));
  nor2 g01787(.a(new_n1980), .b(new_n1978), .O(new_n1981));
  nor2 g01788(.a(new_n1981), .b(new_n1970), .O(new_n1982));
  inv1 g01789(.a(new_n1970), .O(new_n1983));
  inv1 g01790(.a(new_n1981), .O(new_n1984));
  nor2 g01791(.a(new_n1984), .b(new_n1983), .O(new_n1985));
  nor2 g01792(.a(new_n1985), .b(new_n1982), .O(new_n1986));
  inv1 g01793(.a(new_n1986), .O(new_n1987));
  nor2 g01794(.a(new_n1987), .b(new_n1969), .O(new_n1988));
  nor2 g01795(.a(new_n1986), .b(new_n1968), .O(new_n1989));
  nor2 g01796(.a(new_n1989), .b(new_n1988), .O(new_n1990));
  inv1 g01797(.a(new_n1990), .O(new_n1991));
  nor2 g01798(.a(new_n1991), .b(new_n1955), .O(new_n1992));
  nor2 g01799(.a(new_n1990), .b(new_n1954), .O(new_n1993));
  nor2 g01800(.a(new_n1993), .b(new_n1992), .O(new_n1994));
  inv1 g01801(.a(new_n1994), .O(new_n1995));
  nor2 g01802(.a(new_n1995), .b(new_n1901), .O(new_n1996));
  nor2 g01803(.a(new_n1994), .b(new_n1900), .O(new_n1997));
  nor2 g01804(.a(new_n1997), .b(new_n1996), .O(new_n1998));
  nor2 g01805(.a(new_n1998), .b(new_n1869), .O(new_n1999));
  inv1 g01806(.a(new_n1998), .O(new_n2000));
  nor2 g01807(.a(new_n2000), .b(new_n1868), .O(new_n2001));
  nor2 g01808(.a(new_n2001), .b(new_n1999), .O(new_n2002));
  inv1 g01809(.a(new_n2002), .O(new_n2003));
  nor2 g01810(.a(new_n1863), .b(new_n1859), .O(new_n2004));
  nor2 g01811(.a(new_n2004), .b(new_n2003), .O(new_n2005));
  inv1 g01812(.a(new_n2004), .O(new_n2006));
  nor2 g01813(.a(new_n2006), .b(new_n2002), .O(new_n2007));
  nor2 g01814(.a(new_n2007), .b(new_n2005), .O(new_n2008));
  inv1 g01815(.a(new_n2008), .O(\asquared[26] ));
  nor2 g01816(.a(new_n1996), .b(new_n1897), .O(new_n2010));
  nor2 g01817(.a(new_n1992), .b(new_n1951), .O(new_n2011));
  nor2 g01818(.a(new_n1988), .b(new_n1982), .O(new_n2012));
  nor2 g01819(.a(new_n699), .b(new_n569), .O(new_n2013));
  nor2 g01820(.a(new_n1903), .b(new_n194), .O(new_n2014));
  nor2 g01821(.a(new_n2014), .b(new_n2013), .O(new_n2015));
  inv1 g01822(.a(new_n2013), .O(new_n2016));
  inv1 g01823(.a(new_n2014), .O(new_n2017));
  nor2 g01824(.a(new_n2017), .b(new_n2016), .O(new_n2018));
  nor2 g01825(.a(new_n2018), .b(new_n2015), .O(new_n2019));
  inv1 g01826(.a(new_n2019), .O(new_n2020));
  nor2 g01827(.a(new_n1980), .b(new_n1973), .O(new_n2021));
  inv1 g01828(.a(new_n2021), .O(new_n2022));
  nor2 g01829(.a(new_n2022), .b(new_n2020), .O(new_n2023));
  nor2 g01830(.a(new_n2021), .b(new_n2019), .O(new_n2024));
  nor2 g01831(.a(new_n2024), .b(new_n2023), .O(new_n2025));
  inv1 g01832(.a(new_n2025), .O(new_n2026));
  nor2 g01833(.a(new_n1943), .b(new_n1936), .O(new_n2027));
  inv1 g01834(.a(new_n2027), .O(new_n2028));
  nor2 g01835(.a(new_n2028), .b(new_n2026), .O(new_n2029));
  nor2 g01836(.a(new_n2027), .b(new_n2025), .O(new_n2030));
  nor2 g01837(.a(new_n2030), .b(new_n2029), .O(new_n2031));
  inv1 g01838(.a(new_n2031), .O(new_n2032));
  nor2 g01839(.a(new_n1948), .b(new_n1927), .O(new_n2033));
  nor2 g01840(.a(new_n2033), .b(new_n2032), .O(new_n2034));
  inv1 g01841(.a(new_n2033), .O(new_n2035));
  nor2 g01842(.a(new_n2035), .b(new_n2031), .O(new_n2036));
  nor2 g01843(.a(new_n2036), .b(new_n2034), .O(new_n2037));
  inv1 g01844(.a(new_n2037), .O(new_n2038));
  nor2 g01845(.a(new_n2038), .b(new_n2012), .O(new_n2039));
  inv1 g01846(.a(new_n2012), .O(new_n2040));
  nor2 g01847(.a(new_n2037), .b(new_n2040), .O(new_n2041));
  nor2 g01848(.a(new_n2041), .b(new_n2039), .O(new_n2042));
  inv1 g01849(.a(new_n2042), .O(new_n2043));
  nor2 g01850(.a(new_n2043), .b(new_n2011), .O(new_n2044));
  inv1 g01851(.a(new_n2011), .O(new_n2045));
  nor2 g01852(.a(new_n2042), .b(new_n2045), .O(new_n2046));
  nor2 g01853(.a(new_n2046), .b(new_n2044), .O(new_n2047));
  inv1 g01854(.a(new_n2047), .O(new_n2048));
  nor2 g01855(.a(new_n1893), .b(new_n1887), .O(new_n2049));
  inv1 g01856(.a(new_n2049), .O(new_n2050));
  nor2 g01857(.a(new_n1297), .b(new_n257), .O(new_n2051));
  nor2 g01858(.a(new_n1425), .b(new_n229), .O(new_n2052));
  nor2 g01859(.a(new_n2052), .b(new_n2051), .O(new_n2053));
  nor2 g01860(.a(new_n1425), .b(new_n257), .O(new_n2054));
  inv1 g01861(.a(new_n2054), .O(new_n2055));
  nor2 g01862(.a(new_n2055), .b(new_n1605), .O(new_n2056));
  nor2 g01863(.a(new_n2056), .b(new_n2053), .O(new_n2057));
  nor2 g01864(.a(new_n2057), .b(new_n1938), .O(new_n2058));
  inv1 g01865(.a(new_n2057), .O(new_n2059));
  nor2 g01866(.a(new_n2059), .b(new_n1937), .O(new_n2060));
  nor2 g01867(.a(new_n2060), .b(new_n2058), .O(new_n2061));
  nor2 g01868(.a(new_n1736), .b(new_n196), .O(new_n2062));
  inv1 g01869(.a(new_n2062), .O(new_n2063));
  nor2 g01870(.a(new_n1647), .b(new_n203), .O(new_n2064));
  nor2 g01871(.a(new_n1199), .b(new_n295), .O(new_n2065));
  nor2 g01872(.a(new_n2065), .b(new_n2064), .O(new_n2066));
  inv1 g01873(.a(new_n2064), .O(new_n2067));
  inv1 g01874(.a(new_n2065), .O(new_n2068));
  nor2 g01875(.a(new_n2068), .b(new_n2067), .O(new_n2069));
  nor2 g01876(.a(new_n2069), .b(new_n2066), .O(new_n2070));
  nor2 g01877(.a(new_n2070), .b(new_n2063), .O(new_n2071));
  inv1 g01878(.a(new_n2070), .O(new_n2072));
  nor2 g01879(.a(new_n2072), .b(new_n2062), .O(new_n2073));
  nor2 g01880(.a(new_n2073), .b(new_n2071), .O(new_n2074));
  nor2 g01881(.a(new_n847), .b(new_n438), .O(new_n2075));
  nor2 g01882(.a(new_n800), .b(new_n502), .O(new_n2076));
  nor2 g01883(.a(new_n2076), .b(new_n2075), .O(new_n2077));
  nor2 g01884(.a(new_n847), .b(new_n502), .O(new_n2078));
  inv1 g01885(.a(new_n2078), .O(new_n2079));
  nor2 g01886(.a(new_n2079), .b(new_n1780), .O(new_n2080));
  nor2 g01887(.a(new_n2080), .b(new_n2077), .O(new_n2081));
  nor2 g01888(.a(new_n2081), .b(new_n1920), .O(new_n2082));
  inv1 g01889(.a(new_n2081), .O(new_n2083));
  nor2 g01890(.a(new_n2083), .b(new_n1919), .O(new_n2084));
  nor2 g01891(.a(new_n2084), .b(new_n2082), .O(new_n2085));
  nor2 g01892(.a(new_n2085), .b(new_n2074), .O(new_n2086));
  inv1 g01893(.a(new_n2074), .O(new_n2087));
  inv1 g01894(.a(new_n2085), .O(new_n2088));
  nor2 g01895(.a(new_n2088), .b(new_n2087), .O(new_n2089));
  nor2 g01896(.a(new_n2089), .b(new_n2086), .O(new_n2090));
  inv1 g01897(.a(new_n2090), .O(new_n2091));
  nor2 g01898(.a(new_n2091), .b(new_n2061), .O(new_n2092));
  inv1 g01899(.a(new_n2061), .O(new_n2093));
  nor2 g01900(.a(new_n2090), .b(new_n2093), .O(new_n2094));
  nor2 g01901(.a(new_n2094), .b(new_n2092), .O(new_n2095));
  nor2 g01902(.a(new_n2095), .b(new_n2050), .O(new_n2096));
  inv1 g01903(.a(new_n2095), .O(new_n2097));
  nor2 g01904(.a(new_n2097), .b(new_n2049), .O(new_n2098));
  nor2 g01905(.a(new_n2098), .b(new_n2096), .O(new_n2099));
  inv1 g01906(.a(new_n2099), .O(new_n2100));
  nor2 g01907(.a(new_n1881), .b(new_n1875), .O(new_n2101));
  inv1 g01908(.a(new_n2101), .O(new_n2102));
  inv1 g01909(.a(new_n1746), .O(new_n2103));
  nor2 g01910(.a(new_n2103), .b(\a[24] ), .O(new_n2104));
  nor2 g01911(.a(new_n2104), .b(new_n1965), .O(new_n2105));
  inv1 g01912(.a(new_n2105), .O(new_n2106));
  nor2 g01913(.a(new_n2106), .b(new_n2102), .O(new_n2107));
  nor2 g01914(.a(new_n2105), .b(new_n2101), .O(new_n2108));
  nor2 g01915(.a(new_n2108), .b(new_n2107), .O(new_n2109));
  inv1 g01916(.a(new_n2109), .O(new_n2110));
  nor2 g01917(.a(new_n1925), .b(new_n1918), .O(new_n2111));
  nor2 g01918(.a(new_n1912), .b(new_n1905), .O(new_n2112));
  nor2 g01919(.a(new_n2112), .b(new_n2111), .O(new_n2113));
  inv1 g01920(.a(new_n2111), .O(new_n2114));
  inv1 g01921(.a(new_n2112), .O(new_n2115));
  nor2 g01922(.a(new_n2115), .b(new_n2114), .O(new_n2116));
  nor2 g01923(.a(new_n2116), .b(new_n2113), .O(new_n2117));
  inv1 g01924(.a(new_n2117), .O(new_n2118));
  nor2 g01925(.a(new_n1957), .b(new_n613), .O(new_n2119));
  inv1 g01926(.a(new_n2119), .O(new_n2120));
  inv1 g01927(.a(\a[26] ), .O(new_n2121));
  nor2 g01928(.a(new_n2121), .b(new_n198), .O(new_n2122));
  nor2 g01929(.a(new_n1086), .b(new_n322), .O(new_n2123));
  nor2 g01930(.a(new_n2123), .b(new_n2122), .O(new_n2124));
  inv1 g01931(.a(new_n2122), .O(new_n2125));
  inv1 g01932(.a(new_n2123), .O(new_n2126));
  nor2 g01933(.a(new_n2126), .b(new_n2125), .O(new_n2127));
  nor2 g01934(.a(new_n2127), .b(new_n2124), .O(new_n2128));
  nor2 g01935(.a(new_n2128), .b(new_n2120), .O(new_n2129));
  inv1 g01936(.a(new_n2128), .O(new_n2130));
  nor2 g01937(.a(new_n2130), .b(new_n2119), .O(new_n2131));
  nor2 g01938(.a(new_n2131), .b(new_n2129), .O(new_n2132));
  nor2 g01939(.a(new_n2132), .b(new_n2118), .O(new_n2133));
  inv1 g01940(.a(new_n2132), .O(new_n2134));
  nor2 g01941(.a(new_n2134), .b(new_n2117), .O(new_n2135));
  nor2 g01942(.a(new_n2135), .b(new_n2133), .O(new_n2136));
  inv1 g01943(.a(new_n2136), .O(new_n2137));
  nor2 g01944(.a(new_n2137), .b(new_n2110), .O(new_n2138));
  nor2 g01945(.a(new_n2136), .b(new_n2109), .O(new_n2139));
  nor2 g01946(.a(new_n2139), .b(new_n2138), .O(new_n2140));
  inv1 g01947(.a(new_n2140), .O(new_n2141));
  nor2 g01948(.a(new_n2141), .b(new_n2100), .O(new_n2142));
  nor2 g01949(.a(new_n2140), .b(new_n2099), .O(new_n2143));
  nor2 g01950(.a(new_n2143), .b(new_n2142), .O(new_n2144));
  inv1 g01951(.a(new_n2144), .O(new_n2145));
  nor2 g01952(.a(new_n2145), .b(new_n2048), .O(new_n2146));
  nor2 g01953(.a(new_n2144), .b(new_n2047), .O(new_n2147));
  nor2 g01954(.a(new_n2147), .b(new_n2146), .O(new_n2148));
  inv1 g01955(.a(new_n2148), .O(new_n2149));
  nor2 g01956(.a(new_n2149), .b(new_n2010), .O(new_n2150));
  inv1 g01957(.a(new_n2010), .O(new_n2151));
  nor2 g01958(.a(new_n2148), .b(new_n2151), .O(new_n2152));
  nor2 g01959(.a(new_n2152), .b(new_n2150), .O(new_n2153));
  inv1 g01960(.a(new_n2153), .O(new_n2154));
  nor2 g01961(.a(new_n2005), .b(new_n1999), .O(new_n2155));
  nor2 g01962(.a(new_n2155), .b(new_n2154), .O(new_n2156));
  inv1 g01963(.a(new_n2155), .O(new_n2157));
  nor2 g01964(.a(new_n2157), .b(new_n2153), .O(new_n2158));
  nor2 g01965(.a(new_n2158), .b(new_n2156), .O(new_n2159));
  inv1 g01966(.a(new_n2159), .O(\asquared[27] ));
  nor2 g01967(.a(new_n2146), .b(new_n2044), .O(new_n2161));
  nor2 g01968(.a(new_n2142), .b(new_n2098), .O(new_n2162));
  nor2 g01969(.a(new_n2084), .b(new_n2077), .O(new_n2163));
  nor2 g01970(.a(new_n2060), .b(new_n2053), .O(new_n2164));
  nor2 g01971(.a(new_n2164), .b(new_n2163), .O(new_n2165));
  inv1 g01972(.a(new_n2163), .O(new_n2166));
  inv1 g01973(.a(new_n2164), .O(new_n2167));
  nor2 g01974(.a(new_n2167), .b(new_n2166), .O(new_n2168));
  nor2 g01975(.a(new_n2168), .b(new_n2165), .O(new_n2169));
  nor2 g01976(.a(new_n2073), .b(new_n2066), .O(new_n2170));
  nor2 g01977(.a(new_n2170), .b(new_n2169), .O(new_n2171));
  inv1 g01978(.a(new_n2169), .O(new_n2172));
  inv1 g01979(.a(new_n2170), .O(new_n2173));
  nor2 g01980(.a(new_n2173), .b(new_n2172), .O(new_n2174));
  nor2 g01981(.a(new_n2174), .b(new_n2171), .O(new_n2175));
  inv1 g01982(.a(new_n2175), .O(new_n2176));
  nor2 g01983(.a(new_n2138), .b(new_n2108), .O(new_n2177));
  nor2 g01984(.a(new_n2177), .b(new_n2176), .O(new_n2178));
  inv1 g01985(.a(new_n2177), .O(new_n2179));
  nor2 g01986(.a(new_n2179), .b(new_n2175), .O(new_n2180));
  nor2 g01987(.a(new_n2180), .b(new_n2178), .O(new_n2181));
  inv1 g01988(.a(new_n2181), .O(new_n2182));
  inv1 g01989(.a(new_n2018), .O(new_n2183));
  inv1 g01990(.a(\a[27] ), .O(new_n2184));
  nor2 g01991(.a(new_n2184), .b(new_n198), .O(new_n2185));
  inv1 g01992(.a(new_n2185), .O(new_n2186));
  nor2 g01993(.a(new_n2186), .b(new_n2183), .O(new_n2187));
  nor2 g01994(.a(new_n2185), .b(new_n2018), .O(new_n2188));
  nor2 g01995(.a(new_n2188), .b(new_n2187), .O(new_n2189));
  inv1 g01996(.a(new_n2189), .O(new_n2190));
  nor2 g01997(.a(new_n772), .b(new_n2121), .O(new_n2191));
  nor2 g01998(.a(new_n2191), .b(new_n699), .O(new_n2192));
  nor2 g01999(.a(\a[14] ), .b(new_n194), .O(new_n2193));
  inv1 g02000(.a(new_n2193), .O(new_n2194));
  nor2 g02001(.a(new_n2194), .b(new_n2121), .O(new_n2195));
  nor2 g02002(.a(new_n2195), .b(new_n2192), .O(new_n2196));
  nor2 g02003(.a(new_n2196), .b(new_n2190), .O(new_n2197));
  inv1 g02004(.a(new_n2196), .O(new_n2198));
  nor2 g02005(.a(new_n2198), .b(new_n2189), .O(new_n2199));
  nor2 g02006(.a(new_n2199), .b(new_n2197), .O(new_n2200));
  inv1 g02007(.a(new_n2200), .O(new_n2201));
  nor2 g02008(.a(new_n1493), .b(new_n229), .O(new_n2202));
  inv1 g02009(.a(new_n2202), .O(new_n2203));
  nor2 g02010(.a(new_n699), .b(new_n613), .O(new_n2204));
  nor2 g02011(.a(new_n800), .b(new_n569), .O(new_n2205));
  nor2 g02012(.a(new_n2205), .b(new_n2204), .O(new_n2206));
  nor2 g02013(.a(new_n800), .b(new_n613), .O(new_n2207));
  inv1 g02014(.a(new_n2207), .O(new_n2208));
  nor2 g02015(.a(new_n2208), .b(new_n2016), .O(new_n2209));
  nor2 g02016(.a(new_n2209), .b(new_n2206), .O(new_n2210));
  nor2 g02017(.a(new_n2210), .b(new_n2203), .O(new_n2211));
  inv1 g02018(.a(new_n2210), .O(new_n2212));
  nor2 g02019(.a(new_n2212), .b(new_n2202), .O(new_n2213));
  nor2 g02020(.a(new_n2213), .b(new_n2211), .O(new_n2214));
  nor2 g02021(.a(new_n1736), .b(new_n203), .O(new_n2215));
  inv1 g02022(.a(new_n2215), .O(new_n2216));
  nor2 g02023(.a(new_n1647), .b(new_n214), .O(new_n2217));
  nor2 g02024(.a(new_n2217), .b(new_n2054), .O(new_n2218));
  inv1 g02025(.a(new_n2217), .O(new_n2219));
  nor2 g02026(.a(new_n2219), .b(new_n2055), .O(new_n2220));
  nor2 g02027(.a(new_n2220), .b(new_n2218), .O(new_n2221));
  nor2 g02028(.a(new_n2221), .b(new_n2216), .O(new_n2222));
  inv1 g02029(.a(new_n2221), .O(new_n2223));
  nor2 g02030(.a(new_n2223), .b(new_n2215), .O(new_n2224));
  nor2 g02031(.a(new_n2224), .b(new_n2222), .O(new_n2225));
  nor2 g02032(.a(new_n2225), .b(new_n2214), .O(new_n2226));
  inv1 g02033(.a(new_n2214), .O(new_n2227));
  inv1 g02034(.a(new_n2225), .O(new_n2228));
  nor2 g02035(.a(new_n2228), .b(new_n2227), .O(new_n2229));
  nor2 g02036(.a(new_n2229), .b(new_n2226), .O(new_n2230));
  inv1 g02037(.a(new_n2230), .O(new_n2231));
  nor2 g02038(.a(new_n2231), .b(new_n2201), .O(new_n2232));
  nor2 g02039(.a(new_n2230), .b(new_n2200), .O(new_n2233));
  nor2 g02040(.a(new_n2233), .b(new_n2232), .O(new_n2234));
  inv1 g02041(.a(new_n2234), .O(new_n2235));
  nor2 g02042(.a(new_n2235), .b(new_n2182), .O(new_n2236));
  nor2 g02043(.a(new_n2234), .b(new_n2181), .O(new_n2237));
  nor2 g02044(.a(new_n2237), .b(new_n2236), .O(new_n2238));
  inv1 g02045(.a(new_n2238), .O(new_n2239));
  nor2 g02046(.a(new_n2239), .b(new_n2162), .O(new_n2240));
  inv1 g02047(.a(new_n2162), .O(new_n2241));
  nor2 g02048(.a(new_n2238), .b(new_n2241), .O(new_n2242));
  nor2 g02049(.a(new_n2242), .b(new_n2240), .O(new_n2243));
  inv1 g02050(.a(new_n2243), .O(new_n2244));
  nor2 g02051(.a(new_n2039), .b(new_n2034), .O(new_n2245));
  inv1 g02052(.a(new_n2245), .O(new_n2246));
  nor2 g02053(.a(new_n1297), .b(new_n295), .O(new_n2247));
  nor2 g02054(.a(new_n2247), .b(new_n1907), .O(new_n2248));
  nor2 g02055(.a(new_n1903), .b(new_n295), .O(new_n2249));
  inv1 g02056(.a(new_n2249), .O(new_n2250));
  nor2 g02057(.a(new_n2250), .b(new_n1511), .O(new_n2251));
  nor2 g02058(.a(new_n2251), .b(new_n2248), .O(new_n2252));
  nor2 g02059(.a(new_n2252), .b(new_n2078), .O(new_n2253));
  inv1 g02060(.a(new_n2252), .O(new_n2254));
  nor2 g02061(.a(new_n2254), .b(new_n2079), .O(new_n2255));
  nor2 g02062(.a(new_n2255), .b(new_n2253), .O(new_n2256));
  inv1 g02063(.a(new_n2256), .O(new_n2257));
  nor2 g02064(.a(new_n2131), .b(new_n2124), .O(new_n2258));
  inv1 g02065(.a(new_n2258), .O(new_n2259));
  nor2 g02066(.a(new_n2259), .b(new_n2257), .O(new_n2260));
  nor2 g02067(.a(new_n2258), .b(new_n2256), .O(new_n2261));
  nor2 g02068(.a(new_n2261), .b(new_n2260), .O(new_n2262));
  inv1 g02069(.a(new_n2262), .O(new_n2263));
  nor2 g02070(.a(new_n1199), .b(new_n322), .O(new_n2264));
  inv1 g02071(.a(new_n2264), .O(new_n2265));
  nor2 g02072(.a(new_n941), .b(new_n438), .O(new_n2266));
  nor2 g02073(.a(new_n1086), .b(new_n363), .O(new_n2267));
  nor2 g02074(.a(new_n2267), .b(new_n2266), .O(new_n2268));
  nor2 g02075(.a(new_n1086), .b(new_n438), .O(new_n2269));
  inv1 g02076(.a(new_n2269), .O(new_n2270));
  nor2 g02077(.a(new_n2270), .b(new_n1920), .O(new_n2271));
  nor2 g02078(.a(new_n2271), .b(new_n2268), .O(new_n2272));
  nor2 g02079(.a(new_n2272), .b(new_n2265), .O(new_n2273));
  inv1 g02080(.a(new_n2272), .O(new_n2274));
  nor2 g02081(.a(new_n2274), .b(new_n2264), .O(new_n2275));
  nor2 g02082(.a(new_n2275), .b(new_n2273), .O(new_n2276));
  nor2 g02083(.a(new_n2276), .b(new_n2263), .O(new_n2277));
  inv1 g02084(.a(new_n2276), .O(new_n2278));
  nor2 g02085(.a(new_n2278), .b(new_n2262), .O(new_n2279));
  nor2 g02086(.a(new_n2279), .b(new_n2277), .O(new_n2280));
  nor2 g02087(.a(new_n2280), .b(new_n2246), .O(new_n2281));
  inv1 g02088(.a(new_n2280), .O(new_n2282));
  nor2 g02089(.a(new_n2282), .b(new_n2245), .O(new_n2283));
  nor2 g02090(.a(new_n2283), .b(new_n2281), .O(new_n2284));
  inv1 g02091(.a(new_n2284), .O(new_n2285));
  nor2 g02092(.a(new_n2029), .b(new_n2023), .O(new_n2286));
  inv1 g02093(.a(new_n2286), .O(new_n2287));
  nor2 g02094(.a(new_n2133), .b(new_n2116), .O(new_n2288));
  inv1 g02095(.a(new_n2288), .O(new_n2289));
  nor2 g02096(.a(new_n2289), .b(new_n2287), .O(new_n2290));
  nor2 g02097(.a(new_n2288), .b(new_n2286), .O(new_n2291));
  nor2 g02098(.a(new_n2291), .b(new_n2290), .O(new_n2292));
  nor2 g02099(.a(new_n2092), .b(new_n2086), .O(new_n2293));
  inv1 g02100(.a(new_n2293), .O(new_n2294));
  nor2 g02101(.a(new_n2294), .b(new_n2292), .O(new_n2295));
  inv1 g02102(.a(new_n2292), .O(new_n2296));
  nor2 g02103(.a(new_n2293), .b(new_n2296), .O(new_n2297));
  nor2 g02104(.a(new_n2297), .b(new_n2295), .O(new_n2298));
  inv1 g02105(.a(new_n2298), .O(new_n2299));
  nor2 g02106(.a(new_n2299), .b(new_n2285), .O(new_n2300));
  nor2 g02107(.a(new_n2298), .b(new_n2284), .O(new_n2301));
  nor2 g02108(.a(new_n2301), .b(new_n2300), .O(new_n2302));
  inv1 g02109(.a(new_n2302), .O(new_n2303));
  nor2 g02110(.a(new_n2303), .b(new_n2244), .O(new_n2304));
  nor2 g02111(.a(new_n2302), .b(new_n2243), .O(new_n2305));
  nor2 g02112(.a(new_n2305), .b(new_n2304), .O(new_n2306));
  inv1 g02113(.a(new_n2306), .O(new_n2307));
  nor2 g02114(.a(new_n2307), .b(new_n2161), .O(new_n2308));
  inv1 g02115(.a(new_n2161), .O(new_n2309));
  nor2 g02116(.a(new_n2306), .b(new_n2309), .O(new_n2310));
  nor2 g02117(.a(new_n2310), .b(new_n2308), .O(new_n2311));
  inv1 g02118(.a(new_n2311), .O(new_n2312));
  nor2 g02119(.a(new_n2156), .b(new_n2152), .O(new_n2313));
  nor2 g02120(.a(new_n2313), .b(new_n2312), .O(new_n2314));
  inv1 g02121(.a(new_n2313), .O(new_n2315));
  nor2 g02122(.a(new_n2315), .b(new_n2311), .O(new_n2316));
  nor2 g02123(.a(new_n2316), .b(new_n2314), .O(new_n2317));
  inv1 g02124(.a(new_n2317), .O(\asquared[28] ));
  nor2 g02125(.a(new_n2236), .b(new_n2178), .O(new_n2319));
  inv1 g02126(.a(new_n2319), .O(new_n2320));
  nor2 g02127(.a(new_n1425), .b(new_n295), .O(new_n2321));
  inv1 g02128(.a(new_n2321), .O(new_n2322));
  nor2 g02129(.a(new_n1647), .b(new_n229), .O(new_n2323));
  nor2 g02130(.a(new_n2323), .b(new_n1758), .O(new_n2324));
  nor2 g02131(.a(new_n1647), .b(new_n257), .O(new_n2325));
  inv1 g02132(.a(new_n2325), .O(new_n2326));
  nor2 g02133(.a(new_n2326), .b(new_n2203), .O(new_n2327));
  nor2 g02134(.a(new_n2327), .b(new_n2324), .O(new_n2328));
  nor2 g02135(.a(new_n2328), .b(new_n2322), .O(new_n2329));
  inv1 g02136(.a(new_n2328), .O(new_n2330));
  nor2 g02137(.a(new_n2330), .b(new_n2321), .O(new_n2331));
  nor2 g02138(.a(new_n2331), .b(new_n2329), .O(new_n2332));
  nor2 g02139(.a(new_n1297), .b(new_n322), .O(new_n2333));
  inv1 g02140(.a(new_n2333), .O(new_n2334));
  nor2 g02141(.a(new_n1903), .b(new_n203), .O(new_n2335));
  nor2 g02142(.a(new_n1736), .b(new_n214), .O(new_n2336));
  nor2 g02143(.a(new_n2336), .b(new_n2335), .O(new_n2337));
  nor2 g02144(.a(new_n1903), .b(new_n214), .O(new_n2338));
  inv1 g02145(.a(new_n2338), .O(new_n2339));
  nor2 g02146(.a(new_n2339), .b(new_n2216), .O(new_n2340));
  nor2 g02147(.a(new_n2340), .b(new_n2337), .O(new_n2341));
  nor2 g02148(.a(new_n2341), .b(new_n2334), .O(new_n2342));
  inv1 g02149(.a(new_n2341), .O(new_n2343));
  nor2 g02150(.a(new_n2343), .b(new_n2333), .O(new_n2344));
  nor2 g02151(.a(new_n2344), .b(new_n2342), .O(new_n2345));
  nor2 g02152(.a(new_n2197), .b(new_n2187), .O(new_n2346));
  nor2 g02153(.a(new_n2346), .b(new_n2345), .O(new_n2347));
  inv1 g02154(.a(new_n2345), .O(new_n2348));
  inv1 g02155(.a(new_n2346), .O(new_n2349));
  nor2 g02156(.a(new_n2349), .b(new_n2348), .O(new_n2350));
  nor2 g02157(.a(new_n2350), .b(new_n2347), .O(new_n2351));
  inv1 g02158(.a(new_n2351), .O(new_n2352));
  nor2 g02159(.a(new_n2352), .b(new_n2332), .O(new_n2353));
  inv1 g02160(.a(new_n2332), .O(new_n2354));
  nor2 g02161(.a(new_n2351), .b(new_n2354), .O(new_n2355));
  nor2 g02162(.a(new_n2355), .b(new_n2353), .O(new_n2356));
  nor2 g02163(.a(new_n2356), .b(new_n2320), .O(new_n2357));
  inv1 g02164(.a(new_n2356), .O(new_n2358));
  nor2 g02165(.a(new_n2358), .b(new_n2319), .O(new_n2359));
  nor2 g02166(.a(new_n2359), .b(new_n2357), .O(new_n2360));
  inv1 g02167(.a(new_n2360), .O(new_n2361));
  nor2 g02168(.a(new_n2232), .b(new_n2226), .O(new_n2362));
  nor2 g02169(.a(new_n2277), .b(new_n2260), .O(new_n2363));
  inv1 g02170(.a(new_n2191), .O(new_n2364));
  nor2 g02171(.a(new_n2184), .b(new_n194), .O(new_n2365));
  nor2 g02172(.a(new_n2365), .b(new_n2207), .O(new_n2366));
  inv1 g02173(.a(new_n2365), .O(new_n2367));
  nor2 g02174(.a(new_n2367), .b(new_n2208), .O(new_n2368));
  nor2 g02175(.a(new_n2368), .b(new_n2366), .O(new_n2369));
  inv1 g02176(.a(new_n2369), .O(new_n2370));
  nor2 g02177(.a(new_n2370), .b(new_n2364), .O(new_n2371));
  nor2 g02178(.a(new_n2369), .b(new_n2191), .O(new_n2372));
  nor2 g02179(.a(new_n2372), .b(new_n2371), .O(new_n2373));
  inv1 g02180(.a(new_n2373), .O(new_n2374));
  nor2 g02181(.a(new_n2213), .b(new_n2206), .O(new_n2375));
  inv1 g02182(.a(new_n2375), .O(new_n2376));
  nor2 g02183(.a(new_n2376), .b(new_n2374), .O(new_n2377));
  nor2 g02184(.a(new_n2375), .b(new_n2373), .O(new_n2378));
  nor2 g02185(.a(new_n2378), .b(new_n2377), .O(new_n2379));
  inv1 g02186(.a(new_n2379), .O(new_n2380));
  nor2 g02187(.a(new_n2380), .b(new_n2363), .O(new_n2381));
  inv1 g02188(.a(new_n2363), .O(new_n2382));
  nor2 g02189(.a(new_n2379), .b(new_n2382), .O(new_n2383));
  nor2 g02190(.a(new_n2383), .b(new_n2381), .O(new_n2384));
  inv1 g02191(.a(new_n2384), .O(new_n2385));
  nor2 g02192(.a(new_n2385), .b(new_n2362), .O(new_n2386));
  inv1 g02193(.a(new_n2362), .O(new_n2387));
  nor2 g02194(.a(new_n2384), .b(new_n2387), .O(new_n2388));
  nor2 g02195(.a(new_n2388), .b(new_n2386), .O(new_n2389));
  inv1 g02196(.a(new_n2389), .O(new_n2390));
  nor2 g02197(.a(new_n2390), .b(new_n2361), .O(new_n2391));
  nor2 g02198(.a(new_n2389), .b(new_n2360), .O(new_n2392));
  nor2 g02199(.a(new_n2392), .b(new_n2391), .O(new_n2393));
  nor2 g02200(.a(new_n2304), .b(new_n2240), .O(new_n2394));
  nor2 g02201(.a(new_n2300), .b(new_n2283), .O(new_n2395));
  nor2 g02202(.a(new_n2224), .b(new_n2218), .O(new_n2396));
  nor2 g02203(.a(new_n2275), .b(new_n2268), .O(new_n2397));
  nor2 g02204(.a(new_n2397), .b(new_n2396), .O(new_n2398));
  inv1 g02205(.a(new_n2396), .O(new_n2399));
  inv1 g02206(.a(new_n2397), .O(new_n2400));
  nor2 g02207(.a(new_n2400), .b(new_n2399), .O(new_n2401));
  nor2 g02208(.a(new_n2401), .b(new_n2398), .O(new_n2402));
  nor2 g02209(.a(new_n2255), .b(new_n2251), .O(new_n2403));
  inv1 g02210(.a(new_n2403), .O(new_n2404));
  nor2 g02211(.a(new_n2404), .b(new_n2402), .O(new_n2405));
  inv1 g02212(.a(new_n2402), .O(new_n2406));
  nor2 g02213(.a(new_n2403), .b(new_n2406), .O(new_n2407));
  nor2 g02214(.a(new_n2407), .b(new_n2405), .O(new_n2408));
  nor2 g02215(.a(new_n2297), .b(new_n2291), .O(new_n2409));
  inv1 g02216(.a(new_n2409), .O(new_n2410));
  nor2 g02217(.a(new_n2410), .b(new_n2408), .O(new_n2411));
  inv1 g02218(.a(new_n2408), .O(new_n2412));
  nor2 g02219(.a(new_n2409), .b(new_n2412), .O(new_n2413));
  nor2 g02220(.a(new_n2413), .b(new_n2411), .O(new_n2414));
  inv1 g02221(.a(new_n2414), .O(new_n2415));
  nor2 g02222(.a(new_n2174), .b(new_n2168), .O(new_n2416));
  inv1 g02223(.a(new_n2416), .O(new_n2417));
  nor2 g02224(.a(new_n2121), .b(new_n196), .O(new_n2418));
  inv1 g02225(.a(new_n2418), .O(new_n2419));
  nor2 g02226(.a(new_n1199), .b(new_n363), .O(new_n2420));
  nor2 g02227(.a(new_n2420), .b(new_n2269), .O(new_n2421));
  inv1 g02228(.a(new_n2267), .O(new_n2422));
  nor2 g02229(.a(new_n1199), .b(new_n438), .O(new_n2423));
  inv1 g02230(.a(new_n2423), .O(new_n2424));
  nor2 g02231(.a(new_n2424), .b(new_n2422), .O(new_n2425));
  nor2 g02232(.a(new_n2425), .b(new_n2421), .O(new_n2426));
  nor2 g02233(.a(new_n2426), .b(new_n2419), .O(new_n2427));
  inv1 g02234(.a(new_n2426), .O(new_n2428));
  nor2 g02235(.a(new_n2428), .b(new_n2418), .O(new_n2429));
  nor2 g02236(.a(new_n2429), .b(new_n2427), .O(new_n2430));
  nor2 g02237(.a(new_n941), .b(new_n502), .O(new_n2431));
  inv1 g02238(.a(new_n2431), .O(new_n2432));
  inv1 g02239(.a(\a[28] ), .O(new_n2433));
  nor2 g02240(.a(new_n2433), .b(new_n198), .O(new_n2434));
  nor2 g02241(.a(new_n847), .b(new_n569), .O(new_n2435));
  nor2 g02242(.a(new_n2435), .b(new_n2434), .O(new_n2436));
  inv1 g02243(.a(new_n2434), .O(new_n2437));
  inv1 g02244(.a(new_n2435), .O(new_n2438));
  nor2 g02245(.a(new_n2438), .b(new_n2437), .O(new_n2439));
  nor2 g02246(.a(new_n2439), .b(new_n2436), .O(new_n2440));
  nor2 g02247(.a(new_n2440), .b(new_n2432), .O(new_n2441));
  inv1 g02248(.a(new_n2440), .O(new_n2442));
  nor2 g02249(.a(new_n2442), .b(new_n2431), .O(new_n2443));
  nor2 g02250(.a(new_n2443), .b(new_n2441), .O(new_n2444));
  nor2 g02251(.a(new_n2444), .b(new_n2430), .O(new_n2445));
  inv1 g02252(.a(new_n2430), .O(new_n2446));
  inv1 g02253(.a(new_n2444), .O(new_n2447));
  nor2 g02254(.a(new_n2447), .b(new_n2446), .O(new_n2448));
  nor2 g02255(.a(new_n2448), .b(new_n2445), .O(new_n2449));
  nor2 g02256(.a(new_n2449), .b(new_n2417), .O(new_n2450));
  inv1 g02257(.a(new_n2449), .O(new_n2451));
  nor2 g02258(.a(new_n2451), .b(new_n2416), .O(new_n2452));
  nor2 g02259(.a(new_n2452), .b(new_n2450), .O(new_n2453));
  inv1 g02260(.a(new_n2453), .O(new_n2454));
  nor2 g02261(.a(new_n2454), .b(new_n2415), .O(new_n2455));
  nor2 g02262(.a(new_n2453), .b(new_n2414), .O(new_n2456));
  nor2 g02263(.a(new_n2456), .b(new_n2455), .O(new_n2457));
  inv1 g02264(.a(new_n2457), .O(new_n2458));
  nor2 g02265(.a(new_n2458), .b(new_n2395), .O(new_n2459));
  inv1 g02266(.a(new_n2395), .O(new_n2460));
  nor2 g02267(.a(new_n2457), .b(new_n2460), .O(new_n2461));
  nor2 g02268(.a(new_n2461), .b(new_n2459), .O(new_n2462));
  inv1 g02269(.a(new_n2462), .O(new_n2463));
  nor2 g02270(.a(new_n2463), .b(new_n2394), .O(new_n2464));
  inv1 g02271(.a(new_n2394), .O(new_n2465));
  nor2 g02272(.a(new_n2462), .b(new_n2465), .O(new_n2466));
  nor2 g02273(.a(new_n2466), .b(new_n2464), .O(new_n2467));
  nor2 g02274(.a(new_n2467), .b(new_n2393), .O(new_n2468));
  inv1 g02275(.a(new_n2393), .O(new_n2469));
  inv1 g02276(.a(new_n2467), .O(new_n2470));
  nor2 g02277(.a(new_n2470), .b(new_n2469), .O(new_n2471));
  nor2 g02278(.a(new_n2471), .b(new_n2468), .O(new_n2472));
  inv1 g02279(.a(new_n2472), .O(new_n2473));
  nor2 g02280(.a(new_n2314), .b(new_n2310), .O(new_n2474));
  nor2 g02281(.a(new_n2474), .b(new_n2473), .O(new_n2475));
  inv1 g02282(.a(new_n2474), .O(new_n2476));
  nor2 g02283(.a(new_n2476), .b(new_n2472), .O(new_n2477));
  nor2 g02284(.a(new_n2477), .b(new_n2475), .O(new_n2478));
  inv1 g02285(.a(new_n2478), .O(\asquared[29] ));
  nor2 g02286(.a(new_n2464), .b(new_n2459), .O(new_n2480));
  nor2 g02287(.a(new_n2455), .b(new_n2413), .O(new_n2481));
  inv1 g02288(.a(new_n2481), .O(new_n2482));
  nor2 g02289(.a(new_n2386), .b(new_n2381), .O(new_n2483));
  inv1 g02290(.a(new_n2483), .O(new_n2484));
  nor2 g02291(.a(new_n2484), .b(new_n2482), .O(new_n2485));
  nor2 g02292(.a(new_n2483), .b(new_n2481), .O(new_n2486));
  nor2 g02293(.a(new_n2486), .b(new_n2485), .O(new_n2487));
  inv1 g02294(.a(new_n2487), .O(new_n2488));
  nor2 g02295(.a(new_n2452), .b(new_n2445), .O(new_n2489));
  inv1 g02296(.a(new_n2489), .O(new_n2490));
  nor2 g02297(.a(new_n2353), .b(new_n2347), .O(new_n2491));
  inv1 g02298(.a(new_n2491), .O(new_n2492));
  nor2 g02299(.a(new_n2492), .b(new_n2490), .O(new_n2493));
  nor2 g02300(.a(new_n2491), .b(new_n2489), .O(new_n2494));
  nor2 g02301(.a(new_n2494), .b(new_n2493), .O(new_n2495));
  inv1 g02302(.a(new_n2495), .O(new_n2496));
  nor2 g02303(.a(new_n2443), .b(new_n2436), .O(new_n2497));
  nor2 g02304(.a(new_n2429), .b(new_n2421), .O(new_n2498));
  nor2 g02305(.a(new_n2498), .b(new_n2497), .O(new_n2499));
  inv1 g02306(.a(new_n2497), .O(new_n2500));
  inv1 g02307(.a(new_n2498), .O(new_n2501));
  nor2 g02308(.a(new_n2501), .b(new_n2500), .O(new_n2502));
  nor2 g02309(.a(new_n2502), .b(new_n2499), .O(new_n2503));
  inv1 g02310(.a(new_n2503), .O(new_n2504));
  inv1 g02311(.a(new_n2368), .O(new_n2505));
  inv1 g02312(.a(\a[29] ), .O(new_n2506));
  nor2 g02313(.a(new_n2506), .b(new_n198), .O(new_n2507));
  nor2 g02314(.a(new_n2184), .b(new_n196), .O(new_n2508));
  nor2 g02315(.a(new_n2508), .b(new_n2507), .O(new_n2509));
  nor2 g02316(.a(new_n2506), .b(new_n196), .O(new_n2510));
  inv1 g02317(.a(new_n2510), .O(new_n2511));
  nor2 g02318(.a(new_n2511), .b(new_n2186), .O(new_n2512));
  nor2 g02319(.a(new_n2512), .b(new_n2509), .O(new_n2513));
  nor2 g02320(.a(new_n2513), .b(new_n2505), .O(new_n2514));
  inv1 g02321(.a(new_n2513), .O(new_n2515));
  nor2 g02322(.a(new_n2515), .b(new_n2368), .O(new_n2516));
  nor2 g02323(.a(new_n2516), .b(new_n2514), .O(new_n2517));
  nor2 g02324(.a(new_n2517), .b(new_n2504), .O(new_n2518));
  inv1 g02325(.a(new_n2517), .O(new_n2519));
  nor2 g02326(.a(new_n2519), .b(new_n2503), .O(new_n2520));
  nor2 g02327(.a(new_n2520), .b(new_n2518), .O(new_n2521));
  inv1 g02328(.a(new_n2521), .O(new_n2522));
  nor2 g02329(.a(new_n2522), .b(new_n2496), .O(new_n2523));
  nor2 g02330(.a(new_n2521), .b(new_n2495), .O(new_n2524));
  nor2 g02331(.a(new_n2524), .b(new_n2523), .O(new_n2525));
  inv1 g02332(.a(new_n2525), .O(new_n2526));
  nor2 g02333(.a(new_n2526), .b(new_n2488), .O(new_n2527));
  nor2 g02334(.a(new_n2525), .b(new_n2487), .O(new_n2528));
  nor2 g02335(.a(new_n2528), .b(new_n2527), .O(new_n2529));
  inv1 g02336(.a(new_n2529), .O(new_n2530));
  nor2 g02337(.a(new_n2391), .b(new_n2359), .O(new_n2531));
  nor2 g02338(.a(new_n2407), .b(new_n2401), .O(new_n2532));
  inv1 g02339(.a(new_n2532), .O(new_n2533));
  nor2 g02340(.a(new_n2377), .b(new_n2371), .O(new_n2534));
  nor2 g02341(.a(new_n800), .b(new_n699), .O(new_n2535));
  nor2 g02342(.a(new_n847), .b(new_n613), .O(new_n2536));
  nor2 g02343(.a(new_n2536), .b(new_n2535), .O(new_n2537));
  inv1 g02344(.a(new_n2535), .O(new_n2538));
  inv1 g02345(.a(new_n2536), .O(new_n2539));
  nor2 g02346(.a(new_n2539), .b(new_n2538), .O(new_n2540));
  nor2 g02347(.a(new_n2540), .b(new_n2537), .O(new_n2541));
  nor2 g02348(.a(new_n2541), .b(new_n2326), .O(new_n2542));
  inv1 g02349(.a(new_n2541), .O(new_n2543));
  nor2 g02350(.a(new_n2543), .b(new_n2325), .O(new_n2544));
  nor2 g02351(.a(new_n2544), .b(new_n2542), .O(new_n2545));
  nor2 g02352(.a(new_n2545), .b(new_n2534), .O(new_n2546));
  inv1 g02353(.a(new_n2534), .O(new_n2547));
  inv1 g02354(.a(new_n2545), .O(new_n2548));
  nor2 g02355(.a(new_n2548), .b(new_n2547), .O(new_n2549));
  nor2 g02356(.a(new_n2549), .b(new_n2546), .O(new_n2550));
  nor2 g02357(.a(new_n2550), .b(new_n2533), .O(new_n2551));
  inv1 g02358(.a(new_n2550), .O(new_n2552));
  nor2 g02359(.a(new_n2552), .b(new_n2532), .O(new_n2553));
  nor2 g02360(.a(new_n2553), .b(new_n2551), .O(new_n2554));
  inv1 g02361(.a(new_n2554), .O(new_n2555));
  nor2 g02362(.a(new_n871), .b(new_n2433), .O(new_n2556));
  nor2 g02363(.a(new_n2433), .b(new_n194), .O(new_n2557));
  nor2 g02364(.a(new_n2557), .b(\a[15] ), .O(new_n2558));
  nor2 g02365(.a(new_n2558), .b(new_n2556), .O(new_n2559));
  nor2 g02366(.a(new_n2331), .b(new_n2324), .O(new_n2560));
  nor2 g02367(.a(new_n2560), .b(new_n2559), .O(new_n2561));
  inv1 g02368(.a(new_n2559), .O(new_n2562));
  inv1 g02369(.a(new_n2560), .O(new_n2563));
  nor2 g02370(.a(new_n2563), .b(new_n2562), .O(new_n2564));
  nor2 g02371(.a(new_n2564), .b(new_n2561), .O(new_n2565));
  inv1 g02372(.a(new_n2565), .O(new_n2566));
  nor2 g02373(.a(new_n2344), .b(new_n2337), .O(new_n2567));
  inv1 g02374(.a(new_n2567), .O(new_n2568));
  nor2 g02375(.a(new_n2568), .b(new_n2566), .O(new_n2569));
  nor2 g02376(.a(new_n2567), .b(new_n2565), .O(new_n2570));
  nor2 g02377(.a(new_n2570), .b(new_n2569), .O(new_n2571));
  inv1 g02378(.a(new_n2571), .O(new_n2572));
  nor2 g02379(.a(new_n941), .b(new_n569), .O(new_n2573));
  nor2 g02380(.a(new_n2121), .b(new_n203), .O(new_n2574));
  nor2 g02381(.a(new_n1425), .b(new_n322), .O(new_n2575));
  nor2 g02382(.a(new_n2575), .b(new_n2574), .O(new_n2576));
  nor2 g02383(.a(new_n2121), .b(new_n322), .O(new_n2577));
  inv1 g02384(.a(new_n2577), .O(new_n2578));
  nor2 g02385(.a(new_n2578), .b(new_n1788), .O(new_n2579));
  nor2 g02386(.a(new_n2579), .b(new_n2576), .O(new_n2580));
  inv1 g02387(.a(new_n2580), .O(new_n2581));
  nor2 g02388(.a(new_n2581), .b(new_n2573), .O(new_n2582));
  inv1 g02389(.a(new_n2573), .O(new_n2583));
  nor2 g02390(.a(new_n2580), .b(new_n2583), .O(new_n2584));
  nor2 g02391(.a(new_n2584), .b(new_n2582), .O(new_n2585));
  nor2 g02392(.a(new_n1297), .b(new_n363), .O(new_n2586));
  inv1 g02393(.a(new_n2586), .O(new_n2587));
  nor2 g02394(.a(new_n1086), .b(new_n502), .O(new_n2588));
  nor2 g02395(.a(new_n2588), .b(new_n2423), .O(new_n2589));
  nor2 g02396(.a(new_n1199), .b(new_n502), .O(new_n2590));
  inv1 g02397(.a(new_n2590), .O(new_n2591));
  nor2 g02398(.a(new_n2591), .b(new_n2270), .O(new_n2592));
  nor2 g02399(.a(new_n2592), .b(new_n2589), .O(new_n2593));
  nor2 g02400(.a(new_n2593), .b(new_n2587), .O(new_n2594));
  inv1 g02401(.a(new_n2593), .O(new_n2595));
  nor2 g02402(.a(new_n2595), .b(new_n2586), .O(new_n2596));
  nor2 g02403(.a(new_n2596), .b(new_n2594), .O(new_n2597));
  nor2 g02404(.a(new_n2597), .b(new_n2585), .O(new_n2598));
  inv1 g02405(.a(new_n2585), .O(new_n2599));
  inv1 g02406(.a(new_n2597), .O(new_n2600));
  nor2 g02407(.a(new_n2600), .b(new_n2599), .O(new_n2601));
  nor2 g02408(.a(new_n2601), .b(new_n2598), .O(new_n2602));
  inv1 g02409(.a(new_n2602), .O(new_n2603));
  nor2 g02410(.a(new_n1493), .b(new_n295), .O(new_n2604));
  nor2 g02411(.a(new_n1736), .b(new_n229), .O(new_n2605));
  nor2 g02412(.a(new_n2605), .b(new_n2604), .O(new_n2606));
  nor2 g02413(.a(new_n1736), .b(new_n295), .O(new_n2607));
  inv1 g02414(.a(new_n2607), .O(new_n2608));
  nor2 g02415(.a(new_n2608), .b(new_n2203), .O(new_n2609));
  nor2 g02416(.a(new_n2609), .b(new_n2606), .O(new_n2610));
  nor2 g02417(.a(new_n2610), .b(new_n2339), .O(new_n2611));
  inv1 g02418(.a(new_n2610), .O(new_n2612));
  nor2 g02419(.a(new_n2612), .b(new_n2338), .O(new_n2613));
  nor2 g02420(.a(new_n2613), .b(new_n2611), .O(new_n2614));
  nor2 g02421(.a(new_n2614), .b(new_n2603), .O(new_n2615));
  inv1 g02422(.a(new_n2614), .O(new_n2616));
  nor2 g02423(.a(new_n2616), .b(new_n2602), .O(new_n2617));
  nor2 g02424(.a(new_n2617), .b(new_n2615), .O(new_n2618));
  inv1 g02425(.a(new_n2618), .O(new_n2619));
  nor2 g02426(.a(new_n2619), .b(new_n2572), .O(new_n2620));
  nor2 g02427(.a(new_n2618), .b(new_n2571), .O(new_n2621));
  nor2 g02428(.a(new_n2621), .b(new_n2620), .O(new_n2622));
  inv1 g02429(.a(new_n2622), .O(new_n2623));
  nor2 g02430(.a(new_n2623), .b(new_n2555), .O(new_n2624));
  nor2 g02431(.a(new_n2622), .b(new_n2554), .O(new_n2625));
  nor2 g02432(.a(new_n2625), .b(new_n2624), .O(new_n2626));
  inv1 g02433(.a(new_n2626), .O(new_n2627));
  nor2 g02434(.a(new_n2627), .b(new_n2531), .O(new_n2628));
  inv1 g02435(.a(new_n2531), .O(new_n2629));
  nor2 g02436(.a(new_n2626), .b(new_n2629), .O(new_n2630));
  nor2 g02437(.a(new_n2630), .b(new_n2628), .O(new_n2631));
  inv1 g02438(.a(new_n2631), .O(new_n2632));
  nor2 g02439(.a(new_n2632), .b(new_n2530), .O(new_n2633));
  nor2 g02440(.a(new_n2631), .b(new_n2529), .O(new_n2634));
  nor2 g02441(.a(new_n2634), .b(new_n2633), .O(new_n2635));
  inv1 g02442(.a(new_n2635), .O(new_n2636));
  nor2 g02443(.a(new_n2636), .b(new_n2480), .O(new_n2637));
  inv1 g02444(.a(new_n2480), .O(new_n2638));
  nor2 g02445(.a(new_n2635), .b(new_n2638), .O(new_n2639));
  nor2 g02446(.a(new_n2639), .b(new_n2637), .O(new_n2640));
  inv1 g02447(.a(new_n2640), .O(new_n2641));
  nor2 g02448(.a(new_n2475), .b(new_n2468), .O(new_n2642));
  nor2 g02449(.a(new_n2642), .b(new_n2641), .O(new_n2643));
  inv1 g02450(.a(new_n2642), .O(new_n2644));
  nor2 g02451(.a(new_n2644), .b(new_n2640), .O(new_n2645));
  nor2 g02452(.a(new_n2645), .b(new_n2643), .O(new_n2646));
  inv1 g02453(.a(new_n2646), .O(\asquared[30] ));
  nor2 g02454(.a(new_n2633), .b(new_n2628), .O(new_n2648));
  nor2 g02455(.a(new_n2569), .b(new_n2564), .O(new_n2649));
  inv1 g02456(.a(new_n2649), .O(new_n2650));
  nor2 g02457(.a(new_n847), .b(new_n699), .O(new_n2651));
  nor2 g02458(.a(new_n2506), .b(new_n194), .O(new_n2652));
  nor2 g02459(.a(new_n2652), .b(new_n2651), .O(new_n2653));
  inv1 g02460(.a(new_n2651), .O(new_n2654));
  inv1 g02461(.a(new_n2652), .O(new_n2655));
  nor2 g02462(.a(new_n2655), .b(new_n2654), .O(new_n2656));
  nor2 g02463(.a(new_n2656), .b(new_n2653), .O(new_n2657));
  inv1 g02464(.a(new_n2657), .O(new_n2658));
  inv1 g02465(.a(new_n2556), .O(new_n2659));
  inv1 g02466(.a(\a[30] ), .O(new_n2660));
  nor2 g02467(.a(new_n2660), .b(new_n198), .O(new_n2661));
  inv1 g02468(.a(new_n2661), .O(new_n2662));
  nor2 g02469(.a(new_n2662), .b(new_n2659), .O(new_n2663));
  nor2 g02470(.a(new_n2661), .b(new_n2556), .O(new_n2664));
  nor2 g02471(.a(new_n2664), .b(new_n2663), .O(new_n2665));
  inv1 g02472(.a(new_n2665), .O(new_n2666));
  nor2 g02473(.a(new_n2666), .b(new_n2658), .O(new_n2667));
  nor2 g02474(.a(new_n2665), .b(new_n2657), .O(new_n2668));
  nor2 g02475(.a(new_n2668), .b(new_n2667), .O(new_n2669));
  nor2 g02476(.a(new_n2669), .b(new_n2650), .O(new_n2670));
  inv1 g02477(.a(new_n2669), .O(new_n2671));
  nor2 g02478(.a(new_n2671), .b(new_n2649), .O(new_n2672));
  nor2 g02479(.a(new_n2672), .b(new_n2670), .O(new_n2673));
  nor2 g02480(.a(new_n2518), .b(new_n2502), .O(new_n2674));
  inv1 g02481(.a(new_n2674), .O(new_n2675));
  nor2 g02482(.a(new_n2675), .b(new_n2673), .O(new_n2676));
  inv1 g02483(.a(new_n2673), .O(new_n2677));
  nor2 g02484(.a(new_n2674), .b(new_n2677), .O(new_n2678));
  nor2 g02485(.a(new_n2678), .b(new_n2676), .O(new_n2679));
  nor2 g02486(.a(new_n2624), .b(new_n2620), .O(new_n2680));
  inv1 g02487(.a(new_n2680), .O(new_n2681));
  nor2 g02488(.a(new_n2681), .b(new_n2679), .O(new_n2682));
  inv1 g02489(.a(new_n2679), .O(new_n2683));
  nor2 g02490(.a(new_n2680), .b(new_n2683), .O(new_n2684));
  nor2 g02491(.a(new_n2684), .b(new_n2682), .O(new_n2685));
  inv1 g02492(.a(new_n2685), .O(new_n2686));
  nor2 g02493(.a(new_n2615), .b(new_n2598), .O(new_n2687));
  inv1 g02494(.a(new_n2687), .O(new_n2688));
  nor2 g02495(.a(new_n2544), .b(new_n2537), .O(new_n2689));
  nor2 g02496(.a(new_n2613), .b(new_n2606), .O(new_n2690));
  nor2 g02497(.a(new_n2690), .b(new_n2689), .O(new_n2691));
  inv1 g02498(.a(new_n2689), .O(new_n2692));
  inv1 g02499(.a(new_n2690), .O(new_n2693));
  nor2 g02500(.a(new_n2693), .b(new_n2692), .O(new_n2694));
  nor2 g02501(.a(new_n2694), .b(new_n2691), .O(new_n2695));
  inv1 g02502(.a(new_n2695), .O(new_n2696));
  nor2 g02503(.a(new_n941), .b(new_n613), .O(new_n2697));
  inv1 g02504(.a(new_n2697), .O(new_n2698));
  nor2 g02505(.a(new_n2433), .b(new_n196), .O(new_n2699));
  nor2 g02506(.a(new_n1425), .b(new_n363), .O(new_n2700));
  nor2 g02507(.a(new_n2700), .b(new_n2699), .O(new_n2701));
  inv1 g02508(.a(new_n2699), .O(new_n2702));
  inv1 g02509(.a(new_n2700), .O(new_n2703));
  nor2 g02510(.a(new_n2703), .b(new_n2702), .O(new_n2704));
  nor2 g02511(.a(new_n2704), .b(new_n2701), .O(new_n2705));
  nor2 g02512(.a(new_n2705), .b(new_n2698), .O(new_n2706));
  inv1 g02513(.a(new_n2705), .O(new_n2707));
  nor2 g02514(.a(new_n2707), .b(new_n2697), .O(new_n2708));
  nor2 g02515(.a(new_n2708), .b(new_n2706), .O(new_n2709));
  nor2 g02516(.a(new_n2709), .b(new_n2696), .O(new_n2710));
  inv1 g02517(.a(new_n2709), .O(new_n2711));
  nor2 g02518(.a(new_n2711), .b(new_n2695), .O(new_n2712));
  nor2 g02519(.a(new_n2712), .b(new_n2710), .O(new_n2713));
  nor2 g02520(.a(new_n2713), .b(new_n2688), .O(new_n2714));
  inv1 g02521(.a(new_n2713), .O(new_n2715));
  nor2 g02522(.a(new_n2715), .b(new_n2687), .O(new_n2716));
  nor2 g02523(.a(new_n2716), .b(new_n2714), .O(new_n2717));
  inv1 g02524(.a(new_n2717), .O(new_n2718));
  nor2 g02525(.a(new_n2596), .b(new_n2589), .O(new_n2719));
  nor2 g02526(.a(new_n2582), .b(new_n2576), .O(new_n2720));
  nor2 g02527(.a(new_n2720), .b(new_n2719), .O(new_n2721));
  inv1 g02528(.a(new_n2719), .O(new_n2722));
  inv1 g02529(.a(new_n2720), .O(new_n2723));
  nor2 g02530(.a(new_n2723), .b(new_n2722), .O(new_n2724));
  nor2 g02531(.a(new_n2724), .b(new_n2721), .O(new_n2725));
  nor2 g02532(.a(new_n2516), .b(new_n2509), .O(new_n2726));
  nor2 g02533(.a(new_n2726), .b(new_n2725), .O(new_n2727));
  inv1 g02534(.a(new_n2725), .O(new_n2728));
  inv1 g02535(.a(new_n2726), .O(new_n2729));
  nor2 g02536(.a(new_n2729), .b(new_n2728), .O(new_n2730));
  nor2 g02537(.a(new_n2730), .b(new_n2727), .O(new_n2731));
  inv1 g02538(.a(new_n2731), .O(new_n2732));
  nor2 g02539(.a(new_n2732), .b(new_n2718), .O(new_n2733));
  nor2 g02540(.a(new_n2731), .b(new_n2717), .O(new_n2734));
  nor2 g02541(.a(new_n2734), .b(new_n2733), .O(new_n2735));
  inv1 g02542(.a(new_n2735), .O(new_n2736));
  nor2 g02543(.a(new_n2736), .b(new_n2686), .O(new_n2737));
  nor2 g02544(.a(new_n2735), .b(new_n2685), .O(new_n2738));
  nor2 g02545(.a(new_n2738), .b(new_n2737), .O(new_n2739));
  inv1 g02546(.a(new_n2739), .O(new_n2740));
  nor2 g02547(.a(new_n2527), .b(new_n2486), .O(new_n2741));
  nor2 g02548(.a(new_n2553), .b(new_n2546), .O(new_n2742));
  inv1 g02549(.a(new_n2742), .O(new_n2743));
  nor2 g02550(.a(new_n1297), .b(new_n438), .O(new_n2744));
  inv1 g02551(.a(new_n2744), .O(new_n2745));
  nor2 g02552(.a(new_n1086), .b(new_n569), .O(new_n2746));
  nor2 g02553(.a(new_n2746), .b(new_n2590), .O(new_n2747));
  inv1 g02554(.a(new_n2588), .O(new_n2748));
  nor2 g02555(.a(new_n1199), .b(new_n569), .O(new_n2749));
  inv1 g02556(.a(new_n2749), .O(new_n2750));
  nor2 g02557(.a(new_n2750), .b(new_n2748), .O(new_n2751));
  nor2 g02558(.a(new_n2751), .b(new_n2747), .O(new_n2752));
  nor2 g02559(.a(new_n2752), .b(new_n2745), .O(new_n2753));
  inv1 g02560(.a(new_n2752), .O(new_n2754));
  nor2 g02561(.a(new_n2754), .b(new_n2744), .O(new_n2755));
  nor2 g02562(.a(new_n2755), .b(new_n2753), .O(new_n2756));
  inv1 g02563(.a(new_n2756), .O(new_n2757));
  nor2 g02564(.a(new_n1903), .b(new_n229), .O(new_n2758));
  inv1 g02565(.a(new_n2758), .O(new_n2759));
  nor2 g02566(.a(new_n1647), .b(new_n295), .O(new_n2760));
  nor2 g02567(.a(new_n1736), .b(new_n257), .O(new_n2761));
  nor2 g02568(.a(new_n2761), .b(new_n2760), .O(new_n2762));
  nor2 g02569(.a(new_n2608), .b(new_n2326), .O(new_n2763));
  nor2 g02570(.a(new_n2763), .b(new_n2762), .O(new_n2764));
  nor2 g02571(.a(new_n2764), .b(new_n2759), .O(new_n2765));
  inv1 g02572(.a(new_n2764), .O(new_n2766));
  nor2 g02573(.a(new_n2766), .b(new_n2758), .O(new_n2767));
  nor2 g02574(.a(new_n2767), .b(new_n2765), .O(new_n2768));
  nor2 g02575(.a(new_n2184), .b(new_n203), .O(new_n2769));
  inv1 g02576(.a(new_n2769), .O(new_n2770));
  nor2 g02577(.a(new_n2121), .b(new_n214), .O(new_n2771));
  nor2 g02578(.a(new_n1493), .b(new_n322), .O(new_n2772));
  nor2 g02579(.a(new_n2772), .b(new_n2771), .O(new_n2773));
  inv1 g02580(.a(new_n2771), .O(new_n2774));
  inv1 g02581(.a(new_n2772), .O(new_n2775));
  nor2 g02582(.a(new_n2775), .b(new_n2774), .O(new_n2776));
  nor2 g02583(.a(new_n2776), .b(new_n2773), .O(new_n2777));
  nor2 g02584(.a(new_n2777), .b(new_n2770), .O(new_n2778));
  inv1 g02585(.a(new_n2777), .O(new_n2779));
  nor2 g02586(.a(new_n2779), .b(new_n2769), .O(new_n2780));
  nor2 g02587(.a(new_n2780), .b(new_n2778), .O(new_n2781));
  nor2 g02588(.a(new_n2781), .b(new_n2768), .O(new_n2782));
  inv1 g02589(.a(new_n2768), .O(new_n2783));
  inv1 g02590(.a(new_n2781), .O(new_n2784));
  nor2 g02591(.a(new_n2784), .b(new_n2783), .O(new_n2785));
  nor2 g02592(.a(new_n2785), .b(new_n2782), .O(new_n2786));
  nor2 g02593(.a(new_n2786), .b(new_n2757), .O(new_n2787));
  inv1 g02594(.a(new_n2786), .O(new_n2788));
  nor2 g02595(.a(new_n2788), .b(new_n2756), .O(new_n2789));
  nor2 g02596(.a(new_n2789), .b(new_n2787), .O(new_n2790));
  nor2 g02597(.a(new_n2790), .b(new_n2743), .O(new_n2791));
  inv1 g02598(.a(new_n2790), .O(new_n2792));
  nor2 g02599(.a(new_n2792), .b(new_n2742), .O(new_n2793));
  nor2 g02600(.a(new_n2793), .b(new_n2791), .O(new_n2794));
  inv1 g02601(.a(new_n2794), .O(new_n2795));
  nor2 g02602(.a(new_n2523), .b(new_n2494), .O(new_n2796));
  nor2 g02603(.a(new_n2796), .b(new_n2795), .O(new_n2797));
  inv1 g02604(.a(new_n2796), .O(new_n2798));
  nor2 g02605(.a(new_n2798), .b(new_n2794), .O(new_n2799));
  nor2 g02606(.a(new_n2799), .b(new_n2797), .O(new_n2800));
  inv1 g02607(.a(new_n2800), .O(new_n2801));
  nor2 g02608(.a(new_n2801), .b(new_n2741), .O(new_n2802));
  inv1 g02609(.a(new_n2741), .O(new_n2803));
  nor2 g02610(.a(new_n2800), .b(new_n2803), .O(new_n2804));
  nor2 g02611(.a(new_n2804), .b(new_n2802), .O(new_n2805));
  inv1 g02612(.a(new_n2805), .O(new_n2806));
  nor2 g02613(.a(new_n2806), .b(new_n2740), .O(new_n2807));
  nor2 g02614(.a(new_n2805), .b(new_n2739), .O(new_n2808));
  nor2 g02615(.a(new_n2808), .b(new_n2807), .O(new_n2809));
  inv1 g02616(.a(new_n2809), .O(new_n2810));
  nor2 g02617(.a(new_n2810), .b(new_n2648), .O(new_n2811));
  inv1 g02618(.a(new_n2648), .O(new_n2812));
  nor2 g02619(.a(new_n2809), .b(new_n2812), .O(new_n2813));
  nor2 g02620(.a(new_n2813), .b(new_n2811), .O(new_n2814));
  inv1 g02621(.a(new_n2814), .O(new_n2815));
  nor2 g02622(.a(new_n2643), .b(new_n2639), .O(new_n2816));
  nor2 g02623(.a(new_n2816), .b(new_n2815), .O(new_n2817));
  inv1 g02624(.a(new_n2816), .O(new_n2818));
  nor2 g02625(.a(new_n2818), .b(new_n2814), .O(new_n2819));
  nor2 g02626(.a(new_n2819), .b(new_n2817), .O(new_n2820));
  inv1 g02627(.a(new_n2820), .O(\asquared[31] ));
  nor2 g02628(.a(new_n2807), .b(new_n2802), .O(new_n2822));
  nor2 g02629(.a(new_n2737), .b(new_n2684), .O(new_n2823));
  nor2 g02630(.a(new_n2733), .b(new_n2716), .O(new_n2824));
  nor2 g02631(.a(new_n1425), .b(new_n438), .O(new_n2825));
  inv1 g02632(.a(\a[31] ), .O(new_n2826));
  nor2 g02633(.a(new_n2826), .b(new_n198), .O(new_n2827));
  nor2 g02634(.a(new_n1493), .b(new_n363), .O(new_n2828));
  nor2 g02635(.a(new_n2828), .b(new_n2827), .O(new_n2829));
  nor2 g02636(.a(new_n2826), .b(new_n363), .O(new_n2830));
  inv1 g02637(.a(new_n2830), .O(new_n2831));
  nor2 g02638(.a(new_n2831), .b(new_n1504), .O(new_n2832));
  nor2 g02639(.a(new_n2832), .b(new_n2829), .O(new_n2833));
  inv1 g02640(.a(new_n2833), .O(new_n2834));
  nor2 g02641(.a(new_n2834), .b(new_n2825), .O(new_n2835));
  inv1 g02642(.a(new_n2825), .O(new_n2836));
  nor2 g02643(.a(new_n2833), .b(new_n2836), .O(new_n2837));
  nor2 g02644(.a(new_n2837), .b(new_n2835), .O(new_n2838));
  nor2 g02645(.a(new_n2667), .b(new_n2663), .O(new_n2839));
  nor2 g02646(.a(new_n1297), .b(new_n502), .O(new_n2840));
  inv1 g02647(.a(new_n2840), .O(new_n2841));
  nor2 g02648(.a(new_n1086), .b(new_n613), .O(new_n2842));
  nor2 g02649(.a(new_n2842), .b(new_n2749), .O(new_n2843));
  inv1 g02650(.a(new_n2746), .O(new_n2844));
  nor2 g02651(.a(new_n1199), .b(new_n613), .O(new_n2845));
  inv1 g02652(.a(new_n2845), .O(new_n2846));
  nor2 g02653(.a(new_n2846), .b(new_n2844), .O(new_n2847));
  nor2 g02654(.a(new_n2847), .b(new_n2843), .O(new_n2848));
  nor2 g02655(.a(new_n2848), .b(new_n2841), .O(new_n2849));
  inv1 g02656(.a(new_n2848), .O(new_n2850));
  nor2 g02657(.a(new_n2850), .b(new_n2840), .O(new_n2851));
  nor2 g02658(.a(new_n2851), .b(new_n2849), .O(new_n2852));
  nor2 g02659(.a(new_n2852), .b(new_n2839), .O(new_n2853));
  inv1 g02660(.a(new_n2839), .O(new_n2854));
  inv1 g02661(.a(new_n2852), .O(new_n2855));
  nor2 g02662(.a(new_n2855), .b(new_n2854), .O(new_n2856));
  nor2 g02663(.a(new_n2856), .b(new_n2853), .O(new_n2857));
  inv1 g02664(.a(new_n2857), .O(new_n2858));
  nor2 g02665(.a(new_n2858), .b(new_n2838), .O(new_n2859));
  inv1 g02666(.a(new_n2838), .O(new_n2860));
  nor2 g02667(.a(new_n2857), .b(new_n2860), .O(new_n2861));
  nor2 g02668(.a(new_n2861), .b(new_n2859), .O(new_n2862));
  inv1 g02669(.a(new_n2862), .O(new_n2863));
  nor2 g02670(.a(new_n2433), .b(new_n203), .O(new_n2864));
  nor2 g02671(.a(new_n2184), .b(new_n214), .O(new_n2865));
  nor2 g02672(.a(new_n2865), .b(new_n2864), .O(new_n2866));
  nor2 g02673(.a(new_n2433), .b(new_n214), .O(new_n2867));
  inv1 g02674(.a(new_n2867), .O(new_n2868));
  nor2 g02675(.a(new_n2868), .b(new_n2770), .O(new_n2869));
  nor2 g02676(.a(new_n2869), .b(new_n2866), .O(new_n2870));
  nor2 g02677(.a(new_n2870), .b(new_n2511), .O(new_n2871));
  inv1 g02678(.a(new_n2870), .O(new_n2872));
  nor2 g02679(.a(new_n2872), .b(new_n2510), .O(new_n2873));
  nor2 g02680(.a(new_n2873), .b(new_n2871), .O(new_n2874));
  inv1 g02681(.a(new_n2874), .O(new_n2875));
  nor2 g02682(.a(new_n1647), .b(new_n322), .O(new_n2876));
  nor2 g02683(.a(new_n2121), .b(new_n229), .O(new_n2877));
  nor2 g02684(.a(new_n2877), .b(new_n2607), .O(new_n2878));
  inv1 g02685(.a(new_n2605), .O(new_n2879));
  nor2 g02686(.a(new_n2121), .b(new_n295), .O(new_n2880));
  inv1 g02687(.a(new_n2880), .O(new_n2881));
  nor2 g02688(.a(new_n2881), .b(new_n2879), .O(new_n2882));
  nor2 g02689(.a(new_n2882), .b(new_n2878), .O(new_n2883));
  inv1 g02690(.a(new_n2883), .O(new_n2884));
  nor2 g02691(.a(new_n2884), .b(new_n2876), .O(new_n2885));
  inv1 g02692(.a(new_n2876), .O(new_n2886));
  nor2 g02693(.a(new_n2883), .b(new_n2886), .O(new_n2887));
  nor2 g02694(.a(new_n2887), .b(new_n2885), .O(new_n2888));
  nor2 g02695(.a(new_n1903), .b(new_n257), .O(new_n2889));
  inv1 g02696(.a(new_n2889), .O(new_n2890));
  nor2 g02697(.a(new_n847), .b(new_n800), .O(new_n2891));
  nor2 g02698(.a(new_n941), .b(new_n699), .O(new_n2892));
  nor2 g02699(.a(new_n2892), .b(new_n2891), .O(new_n2893));
  nor2 g02700(.a(new_n941), .b(new_n800), .O(new_n2894));
  inv1 g02701(.a(new_n2894), .O(new_n2895));
  nor2 g02702(.a(new_n2895), .b(new_n2654), .O(new_n2896));
  nor2 g02703(.a(new_n2896), .b(new_n2893), .O(new_n2897));
  nor2 g02704(.a(new_n2897), .b(new_n2890), .O(new_n2898));
  inv1 g02705(.a(new_n2897), .O(new_n2899));
  nor2 g02706(.a(new_n2899), .b(new_n2889), .O(new_n2900));
  nor2 g02707(.a(new_n2900), .b(new_n2898), .O(new_n2901));
  nor2 g02708(.a(new_n2901), .b(new_n2888), .O(new_n2902));
  inv1 g02709(.a(new_n2888), .O(new_n2903));
  inv1 g02710(.a(new_n2901), .O(new_n2904));
  nor2 g02711(.a(new_n2904), .b(new_n2903), .O(new_n2905));
  nor2 g02712(.a(new_n2905), .b(new_n2902), .O(new_n2906));
  nor2 g02713(.a(new_n2906), .b(new_n2875), .O(new_n2907));
  inv1 g02714(.a(new_n2906), .O(new_n2908));
  nor2 g02715(.a(new_n2908), .b(new_n2874), .O(new_n2909));
  nor2 g02716(.a(new_n2909), .b(new_n2907), .O(new_n2910));
  inv1 g02717(.a(new_n2910), .O(new_n2911));
  nor2 g02718(.a(new_n2911), .b(new_n2863), .O(new_n2912));
  nor2 g02719(.a(new_n2910), .b(new_n2862), .O(new_n2913));
  nor2 g02720(.a(new_n2913), .b(new_n2912), .O(new_n2914));
  inv1 g02721(.a(new_n2914), .O(new_n2915));
  nor2 g02722(.a(new_n2915), .b(new_n2824), .O(new_n2916));
  inv1 g02723(.a(new_n2824), .O(new_n2917));
  nor2 g02724(.a(new_n2914), .b(new_n2917), .O(new_n2918));
  nor2 g02725(.a(new_n2918), .b(new_n2916), .O(new_n2919));
  inv1 g02726(.a(new_n2919), .O(new_n2920));
  nor2 g02727(.a(new_n2920), .b(new_n2823), .O(new_n2921));
  inv1 g02728(.a(new_n2823), .O(new_n2922));
  nor2 g02729(.a(new_n2919), .b(new_n2922), .O(new_n2923));
  nor2 g02730(.a(new_n2923), .b(new_n2921), .O(new_n2924));
  inv1 g02731(.a(new_n2924), .O(new_n2925));
  nor2 g02732(.a(new_n2797), .b(new_n2793), .O(new_n2926));
  inv1 g02733(.a(new_n2926), .O(new_n2927));
  nor2 g02734(.a(new_n2730), .b(new_n2724), .O(new_n2928));
  inv1 g02735(.a(new_n2928), .O(new_n2929));
  nor2 g02736(.a(new_n2710), .b(new_n2694), .O(new_n2930));
  inv1 g02737(.a(new_n2930), .O(new_n2931));
  nor2 g02738(.a(new_n2931), .b(new_n2929), .O(new_n2932));
  nor2 g02739(.a(new_n2930), .b(new_n2928), .O(new_n2933));
  nor2 g02740(.a(new_n2933), .b(new_n2932), .O(new_n2934));
  inv1 g02741(.a(new_n2934), .O(new_n2935));
  nor2 g02742(.a(new_n2660), .b(new_n194), .O(new_n2936));
  inv1 g02743(.a(new_n2936), .O(new_n2937));
  nor2 g02744(.a(new_n2656), .b(new_n847), .O(new_n2938));
  nor2 g02745(.a(new_n2938), .b(new_n2937), .O(new_n2939));
  inv1 g02746(.a(new_n2938), .O(new_n2940));
  nor2 g02747(.a(new_n2940), .b(new_n2936), .O(new_n2941));
  nor2 g02748(.a(new_n2941), .b(new_n2939), .O(new_n2942));
  nor2 g02749(.a(new_n2767), .b(new_n2762), .O(new_n2943));
  inv1 g02750(.a(new_n2943), .O(new_n2944));
  nor2 g02751(.a(new_n2944), .b(new_n2942), .O(new_n2945));
  inv1 g02752(.a(new_n2942), .O(new_n2946));
  nor2 g02753(.a(new_n2943), .b(new_n2946), .O(new_n2947));
  nor2 g02754(.a(new_n2947), .b(new_n2945), .O(new_n2948));
  inv1 g02755(.a(new_n2948), .O(new_n2949));
  nor2 g02756(.a(new_n2949), .b(new_n2935), .O(new_n2950));
  nor2 g02757(.a(new_n2948), .b(new_n2934), .O(new_n2951));
  nor2 g02758(.a(new_n2951), .b(new_n2950), .O(new_n2952));
  nor2 g02759(.a(new_n2952), .b(new_n2927), .O(new_n2953));
  inv1 g02760(.a(new_n2952), .O(new_n2954));
  nor2 g02761(.a(new_n2954), .b(new_n2926), .O(new_n2955));
  nor2 g02762(.a(new_n2955), .b(new_n2953), .O(new_n2956));
  inv1 g02763(.a(new_n2956), .O(new_n2957));
  nor2 g02764(.a(new_n2708), .b(new_n2701), .O(new_n2958));
  nor2 g02765(.a(new_n2780), .b(new_n2773), .O(new_n2959));
  nor2 g02766(.a(new_n2959), .b(new_n2958), .O(new_n2960));
  inv1 g02767(.a(new_n2958), .O(new_n2961));
  inv1 g02768(.a(new_n2959), .O(new_n2962));
  nor2 g02769(.a(new_n2962), .b(new_n2961), .O(new_n2963));
  nor2 g02770(.a(new_n2963), .b(new_n2960), .O(new_n2964));
  nor2 g02771(.a(new_n2755), .b(new_n2747), .O(new_n2965));
  nor2 g02772(.a(new_n2965), .b(new_n2964), .O(new_n2966));
  inv1 g02773(.a(new_n2964), .O(new_n2967));
  inv1 g02774(.a(new_n2965), .O(new_n2968));
  nor2 g02775(.a(new_n2968), .b(new_n2967), .O(new_n2969));
  nor2 g02776(.a(new_n2969), .b(new_n2966), .O(new_n2970));
  nor2 g02777(.a(new_n2789), .b(new_n2782), .O(new_n2971));
  inv1 g02778(.a(new_n2971), .O(new_n2972));
  nor2 g02779(.a(new_n2972), .b(new_n2970), .O(new_n2973));
  inv1 g02780(.a(new_n2970), .O(new_n2974));
  nor2 g02781(.a(new_n2971), .b(new_n2974), .O(new_n2975));
  nor2 g02782(.a(new_n2975), .b(new_n2973), .O(new_n2976));
  nor2 g02783(.a(new_n2678), .b(new_n2672), .O(new_n2977));
  inv1 g02784(.a(new_n2977), .O(new_n2978));
  nor2 g02785(.a(new_n2978), .b(new_n2976), .O(new_n2979));
  inv1 g02786(.a(new_n2976), .O(new_n2980));
  nor2 g02787(.a(new_n2977), .b(new_n2980), .O(new_n2981));
  nor2 g02788(.a(new_n2981), .b(new_n2979), .O(new_n2982));
  inv1 g02789(.a(new_n2982), .O(new_n2983));
  nor2 g02790(.a(new_n2983), .b(new_n2957), .O(new_n2984));
  nor2 g02791(.a(new_n2982), .b(new_n2956), .O(new_n2985));
  nor2 g02792(.a(new_n2985), .b(new_n2984), .O(new_n2986));
  inv1 g02793(.a(new_n2986), .O(new_n2987));
  nor2 g02794(.a(new_n2987), .b(new_n2925), .O(new_n2988));
  nor2 g02795(.a(new_n2986), .b(new_n2924), .O(new_n2989));
  nor2 g02796(.a(new_n2989), .b(new_n2988), .O(new_n2990));
  inv1 g02797(.a(new_n2990), .O(new_n2991));
  nor2 g02798(.a(new_n2991), .b(new_n2822), .O(new_n2992));
  inv1 g02799(.a(new_n2822), .O(new_n2993));
  nor2 g02800(.a(new_n2990), .b(new_n2993), .O(new_n2994));
  nor2 g02801(.a(new_n2994), .b(new_n2992), .O(new_n2995));
  inv1 g02802(.a(new_n2995), .O(new_n2996));
  nor2 g02803(.a(new_n2817), .b(new_n2813), .O(new_n2997));
  nor2 g02804(.a(new_n2997), .b(new_n2996), .O(new_n2998));
  inv1 g02805(.a(new_n2997), .O(new_n2999));
  nor2 g02806(.a(new_n2999), .b(new_n2995), .O(new_n3000));
  nor2 g02807(.a(new_n3000), .b(new_n2998), .O(new_n3001));
  inv1 g02808(.a(new_n3001), .O(\asquared[32] ));
  nor2 g02809(.a(new_n2988), .b(new_n2921), .O(new_n3003));
  nor2 g02810(.a(new_n2984), .b(new_n2955), .O(new_n3004));
  nor2 g02811(.a(new_n2981), .b(new_n2975), .O(new_n3005));
  inv1 g02812(.a(new_n2656), .O(new_n3006));
  nor2 g02813(.a(new_n3006), .b(\a[30] ), .O(new_n3007));
  nor2 g02814(.a(new_n3007), .b(new_n2945), .O(new_n3008));
  inv1 g02815(.a(new_n3008), .O(new_n3009));
  nor2 g02816(.a(new_n1647), .b(new_n363), .O(new_n3010));
  nor2 g02817(.a(new_n2184), .b(new_n229), .O(new_n3011));
  nor2 g02818(.a(new_n3011), .b(new_n2867), .O(new_n3012));
  inv1 g02819(.a(new_n2865), .O(new_n3013));
  nor2 g02820(.a(new_n2433), .b(new_n229), .O(new_n3014));
  inv1 g02821(.a(new_n3014), .O(new_n3015));
  nor2 g02822(.a(new_n3015), .b(new_n3013), .O(new_n3016));
  nor2 g02823(.a(new_n3016), .b(new_n3012), .O(new_n3017));
  inv1 g02824(.a(new_n3017), .O(new_n3018));
  nor2 g02825(.a(new_n3018), .b(new_n3010), .O(new_n3019));
  inv1 g02826(.a(new_n3010), .O(new_n3020));
  nor2 g02827(.a(new_n3017), .b(new_n3020), .O(new_n3021));
  nor2 g02828(.a(new_n3021), .b(new_n3019), .O(new_n3022));
  nor2 g02829(.a(new_n1736), .b(new_n322), .O(new_n3023));
  inv1 g02830(.a(new_n3023), .O(new_n3024));
  nor2 g02831(.a(new_n2121), .b(new_n257), .O(new_n3025));
  nor2 g02832(.a(new_n3025), .b(new_n2249), .O(new_n3026));
  nor2 g02833(.a(new_n2890), .b(new_n2881), .O(new_n3027));
  nor2 g02834(.a(new_n3027), .b(new_n3026), .O(new_n3028));
  nor2 g02835(.a(new_n3028), .b(new_n3024), .O(new_n3029));
  inv1 g02836(.a(new_n3028), .O(new_n3030));
  nor2 g02837(.a(new_n3030), .b(new_n3023), .O(new_n3031));
  nor2 g02838(.a(new_n3031), .b(new_n3029), .O(new_n3032));
  nor2 g02839(.a(new_n3032), .b(new_n3022), .O(new_n3033));
  inv1 g02840(.a(new_n3022), .O(new_n3034));
  inv1 g02841(.a(new_n3032), .O(new_n3035));
  nor2 g02842(.a(new_n3035), .b(new_n3034), .O(new_n3036));
  nor2 g02843(.a(new_n3036), .b(new_n3033), .O(new_n3037));
  nor2 g02844(.a(new_n3037), .b(new_n3009), .O(new_n3038));
  inv1 g02845(.a(new_n3037), .O(new_n3039));
  nor2 g02846(.a(new_n3039), .b(new_n3008), .O(new_n3040));
  nor2 g02847(.a(new_n3040), .b(new_n3038), .O(new_n3041));
  nor2 g02848(.a(new_n1086), .b(new_n699), .O(new_n3042));
  inv1 g02849(.a(new_n3042), .O(new_n3043));
  nor2 g02850(.a(new_n2506), .b(new_n203), .O(new_n3044));
  nor2 g02851(.a(new_n1493), .b(new_n438), .O(new_n3045));
  nor2 g02852(.a(new_n3045), .b(new_n3044), .O(new_n3046));
  inv1 g02853(.a(new_n3044), .O(new_n3047));
  inv1 g02854(.a(new_n3045), .O(new_n3048));
  nor2 g02855(.a(new_n3048), .b(new_n3047), .O(new_n3049));
  nor2 g02856(.a(new_n3049), .b(new_n3046), .O(new_n3050));
  nor2 g02857(.a(new_n3050), .b(new_n3043), .O(new_n3051));
  inv1 g02858(.a(new_n3050), .O(new_n3052));
  nor2 g02859(.a(new_n3052), .b(new_n3042), .O(new_n3053));
  nor2 g02860(.a(new_n3053), .b(new_n3051), .O(new_n3054));
  inv1 g02861(.a(new_n3054), .O(new_n3055));
  nor2 g02862(.a(new_n2937), .b(new_n847), .O(new_n3056));
  inv1 g02863(.a(\a[32] ), .O(new_n3057));
  nor2 g02864(.a(new_n3057), .b(new_n198), .O(new_n3058));
  nor2 g02865(.a(new_n2660), .b(new_n196), .O(new_n3059));
  nor2 g02866(.a(new_n3059), .b(new_n3058), .O(new_n3060));
  nor2 g02867(.a(new_n3057), .b(new_n196), .O(new_n3061));
  inv1 g02868(.a(new_n3061), .O(new_n3062));
  nor2 g02869(.a(new_n3062), .b(new_n2662), .O(new_n3063));
  nor2 g02870(.a(new_n3063), .b(new_n3060), .O(new_n3064));
  inv1 g02871(.a(new_n3064), .O(new_n3065));
  nor2 g02872(.a(new_n3065), .b(new_n3056), .O(new_n3066));
  inv1 g02873(.a(new_n3056), .O(new_n3067));
  nor2 g02874(.a(new_n3064), .b(new_n3067), .O(new_n3068));
  nor2 g02875(.a(new_n3068), .b(new_n3066), .O(new_n3069));
  nor2 g02876(.a(new_n1425), .b(new_n502), .O(new_n3070));
  inv1 g02877(.a(new_n3070), .O(new_n3071));
  nor2 g02878(.a(new_n1297), .b(new_n569), .O(new_n3072));
  nor2 g02879(.a(new_n3072), .b(new_n2845), .O(new_n3073));
  nor2 g02880(.a(new_n1297), .b(new_n613), .O(new_n3074));
  inv1 g02881(.a(new_n3074), .O(new_n3075));
  nor2 g02882(.a(new_n3075), .b(new_n2750), .O(new_n3076));
  nor2 g02883(.a(new_n3076), .b(new_n3073), .O(new_n3077));
  nor2 g02884(.a(new_n3077), .b(new_n3071), .O(new_n3078));
  inv1 g02885(.a(new_n3077), .O(new_n3079));
  nor2 g02886(.a(new_n3079), .b(new_n3070), .O(new_n3080));
  nor2 g02887(.a(new_n3080), .b(new_n3078), .O(new_n3081));
  nor2 g02888(.a(new_n3081), .b(new_n3069), .O(new_n3082));
  inv1 g02889(.a(new_n3069), .O(new_n3083));
  inv1 g02890(.a(new_n3081), .O(new_n3084));
  nor2 g02891(.a(new_n3084), .b(new_n3083), .O(new_n3085));
  nor2 g02892(.a(new_n3085), .b(new_n3082), .O(new_n3086));
  nor2 g02893(.a(new_n3086), .b(new_n3055), .O(new_n3087));
  inv1 g02894(.a(new_n3086), .O(new_n3088));
  nor2 g02895(.a(new_n3088), .b(new_n3054), .O(new_n3089));
  nor2 g02896(.a(new_n3089), .b(new_n3087), .O(new_n3090));
  nor2 g02897(.a(new_n3090), .b(new_n3041), .O(new_n3091));
  inv1 g02898(.a(new_n3041), .O(new_n3092));
  inv1 g02899(.a(new_n3090), .O(new_n3093));
  nor2 g02900(.a(new_n3093), .b(new_n3092), .O(new_n3094));
  nor2 g02901(.a(new_n3094), .b(new_n3091), .O(new_n3095));
  inv1 g02902(.a(new_n3095), .O(new_n3096));
  nor2 g02903(.a(new_n3096), .b(new_n3005), .O(new_n3097));
  inv1 g02904(.a(new_n3005), .O(new_n3098));
  nor2 g02905(.a(new_n3095), .b(new_n3098), .O(new_n3099));
  nor2 g02906(.a(new_n3099), .b(new_n3097), .O(new_n3100));
  inv1 g02907(.a(new_n3100), .O(new_n3101));
  nor2 g02908(.a(new_n3101), .b(new_n3004), .O(new_n3102));
  inv1 g02909(.a(new_n3004), .O(new_n3103));
  nor2 g02910(.a(new_n3100), .b(new_n3103), .O(new_n3104));
  nor2 g02911(.a(new_n3104), .b(new_n3102), .O(new_n3105));
  inv1 g02912(.a(new_n3105), .O(new_n3106));
  nor2 g02913(.a(new_n2950), .b(new_n2933), .O(new_n3107));
  inv1 g02914(.a(new_n3107), .O(new_n3108));
  nor2 g02915(.a(new_n2851), .b(new_n2843), .O(new_n3109));
  nor2 g02916(.a(new_n2835), .b(new_n2829), .O(new_n3110));
  nor2 g02917(.a(new_n3110), .b(new_n3109), .O(new_n3111));
  inv1 g02918(.a(new_n3109), .O(new_n3112));
  inv1 g02919(.a(new_n3110), .O(new_n3113));
  nor2 g02920(.a(new_n3113), .b(new_n3112), .O(new_n3114));
  nor2 g02921(.a(new_n3114), .b(new_n3111), .O(new_n3115));
  nor2 g02922(.a(new_n2873), .b(new_n2866), .O(new_n3116));
  nor2 g02923(.a(new_n3116), .b(new_n3115), .O(new_n3117));
  inv1 g02924(.a(new_n3115), .O(new_n3118));
  inv1 g02925(.a(new_n3116), .O(new_n3119));
  nor2 g02926(.a(new_n3119), .b(new_n3118), .O(new_n3120));
  nor2 g02927(.a(new_n3120), .b(new_n3117), .O(new_n3121));
  inv1 g02928(.a(new_n3121), .O(new_n3122));
  nor2 g02929(.a(new_n2826), .b(new_n194), .O(new_n3123));
  nor2 g02930(.a(new_n3123), .b(new_n2894), .O(new_n3124));
  inv1 g02931(.a(new_n3123), .O(new_n3125));
  nor2 g02932(.a(new_n3125), .b(new_n2895), .O(new_n3126));
  nor2 g02933(.a(new_n3126), .b(new_n3124), .O(new_n3127));
  nor2 g02934(.a(new_n2900), .b(new_n2893), .O(new_n3128));
  nor2 g02935(.a(new_n3128), .b(new_n3127), .O(new_n3129));
  inv1 g02936(.a(new_n3127), .O(new_n3130));
  inv1 g02937(.a(new_n3128), .O(new_n3131));
  nor2 g02938(.a(new_n3131), .b(new_n3130), .O(new_n3132));
  nor2 g02939(.a(new_n3132), .b(new_n3129), .O(new_n3133));
  inv1 g02940(.a(new_n3133), .O(new_n3134));
  nor2 g02941(.a(new_n2885), .b(new_n2878), .O(new_n3135));
  inv1 g02942(.a(new_n3135), .O(new_n3136));
  nor2 g02943(.a(new_n3136), .b(new_n3134), .O(new_n3137));
  nor2 g02944(.a(new_n3135), .b(new_n3133), .O(new_n3138));
  nor2 g02945(.a(new_n3138), .b(new_n3137), .O(new_n3139));
  inv1 g02946(.a(new_n3139), .O(new_n3140));
  nor2 g02947(.a(new_n3140), .b(new_n3122), .O(new_n3141));
  nor2 g02948(.a(new_n3139), .b(new_n3121), .O(new_n3142));
  nor2 g02949(.a(new_n3142), .b(new_n3141), .O(new_n3143));
  nor2 g02950(.a(new_n3143), .b(new_n3108), .O(new_n3144));
  inv1 g02951(.a(new_n3143), .O(new_n3145));
  nor2 g02952(.a(new_n3145), .b(new_n3107), .O(new_n3146));
  nor2 g02953(.a(new_n3146), .b(new_n3144), .O(new_n3147));
  inv1 g02954(.a(new_n3147), .O(new_n3148));
  nor2 g02955(.a(new_n2859), .b(new_n2853), .O(new_n3149));
  inv1 g02956(.a(new_n3149), .O(new_n3150));
  nor2 g02957(.a(new_n2969), .b(new_n2963), .O(new_n3151));
  inv1 g02958(.a(new_n3151), .O(new_n3152));
  nor2 g02959(.a(new_n3152), .b(new_n3150), .O(new_n3153));
  nor2 g02960(.a(new_n3151), .b(new_n3149), .O(new_n3154));
  nor2 g02961(.a(new_n3154), .b(new_n3153), .O(new_n3155));
  nor2 g02962(.a(new_n2909), .b(new_n2902), .O(new_n3156));
  inv1 g02963(.a(new_n3156), .O(new_n3157));
  nor2 g02964(.a(new_n3157), .b(new_n3155), .O(new_n3158));
  inv1 g02965(.a(new_n3155), .O(new_n3159));
  nor2 g02966(.a(new_n3156), .b(new_n3159), .O(new_n3160));
  nor2 g02967(.a(new_n3160), .b(new_n3158), .O(new_n3161));
  nor2 g02968(.a(new_n2916), .b(new_n2912), .O(new_n3162));
  inv1 g02969(.a(new_n3162), .O(new_n3163));
  nor2 g02970(.a(new_n3163), .b(new_n3161), .O(new_n3164));
  inv1 g02971(.a(new_n3161), .O(new_n3165));
  nor2 g02972(.a(new_n3162), .b(new_n3165), .O(new_n3166));
  nor2 g02973(.a(new_n3166), .b(new_n3164), .O(new_n3167));
  inv1 g02974(.a(new_n3167), .O(new_n3168));
  nor2 g02975(.a(new_n3168), .b(new_n3148), .O(new_n3169));
  nor2 g02976(.a(new_n3167), .b(new_n3147), .O(new_n3170));
  nor2 g02977(.a(new_n3170), .b(new_n3169), .O(new_n3171));
  inv1 g02978(.a(new_n3171), .O(new_n3172));
  nor2 g02979(.a(new_n3172), .b(new_n3106), .O(new_n3173));
  nor2 g02980(.a(new_n3171), .b(new_n3105), .O(new_n3174));
  nor2 g02981(.a(new_n3174), .b(new_n3173), .O(new_n3175));
  inv1 g02982(.a(new_n3175), .O(new_n3176));
  nor2 g02983(.a(new_n3176), .b(new_n3003), .O(new_n3177));
  inv1 g02984(.a(new_n3003), .O(new_n3178));
  nor2 g02985(.a(new_n3175), .b(new_n3178), .O(new_n3179));
  nor2 g02986(.a(new_n3179), .b(new_n3177), .O(new_n3180));
  inv1 g02987(.a(new_n3180), .O(new_n3181));
  nor2 g02988(.a(new_n2998), .b(new_n2994), .O(new_n3182));
  nor2 g02989(.a(new_n3182), .b(new_n3181), .O(new_n3183));
  inv1 g02990(.a(new_n3182), .O(new_n3184));
  nor2 g02991(.a(new_n3184), .b(new_n3180), .O(new_n3185));
  nor2 g02992(.a(new_n3185), .b(new_n3183), .O(new_n3186));
  inv1 g02993(.a(new_n3186), .O(\asquared[33] ));
  nor2 g02994(.a(new_n3120), .b(new_n3114), .O(new_n3188));
  inv1 g02995(.a(new_n3188), .O(new_n3189));
  nor2 g02996(.a(new_n3089), .b(new_n3082), .O(new_n3190));
  inv1 g02997(.a(new_n3190), .O(new_n3191));
  nor2 g02998(.a(new_n3191), .b(new_n3189), .O(new_n3192));
  nor2 g02999(.a(new_n3190), .b(new_n3188), .O(new_n3193));
  nor2 g03000(.a(new_n3193), .b(new_n3192), .O(new_n3194));
  nor2 g03001(.a(new_n3040), .b(new_n3033), .O(new_n3195));
  inv1 g03002(.a(new_n3195), .O(new_n3196));
  nor2 g03003(.a(new_n3196), .b(new_n3194), .O(new_n3197));
  inv1 g03004(.a(new_n3194), .O(new_n3198));
  nor2 g03005(.a(new_n3195), .b(new_n3198), .O(new_n3199));
  nor2 g03006(.a(new_n3199), .b(new_n3197), .O(new_n3200));
  inv1 g03007(.a(new_n3200), .O(new_n3201));
  nor2 g03008(.a(new_n3097), .b(new_n3094), .O(new_n3202));
  nor2 g03009(.a(new_n3202), .b(new_n3201), .O(new_n3203));
  inv1 g03010(.a(new_n3202), .O(new_n3204));
  nor2 g03011(.a(new_n3204), .b(new_n3200), .O(new_n3205));
  nor2 g03012(.a(new_n3205), .b(new_n3203), .O(new_n3206));
  inv1 g03013(.a(new_n3206), .O(new_n3207));
  nor2 g03014(.a(new_n3080), .b(new_n3073), .O(new_n3208));
  nor2 g03015(.a(new_n3066), .b(new_n3060), .O(new_n3209));
  nor2 g03016(.a(new_n3209), .b(new_n3208), .O(new_n3210));
  inv1 g03017(.a(new_n3208), .O(new_n3211));
  inv1 g03018(.a(new_n3209), .O(new_n3212));
  nor2 g03019(.a(new_n3212), .b(new_n3211), .O(new_n3213));
  nor2 g03020(.a(new_n3213), .b(new_n3210), .O(new_n3214));
  nor2 g03021(.a(new_n3053), .b(new_n3046), .O(new_n3215));
  nor2 g03022(.a(new_n3215), .b(new_n3214), .O(new_n3216));
  inv1 g03023(.a(new_n3214), .O(new_n3217));
  inv1 g03024(.a(new_n3215), .O(new_n3218));
  nor2 g03025(.a(new_n3218), .b(new_n3217), .O(new_n3219));
  nor2 g03026(.a(new_n3219), .b(new_n3216), .O(new_n3220));
  nor2 g03027(.a(new_n3031), .b(new_n3026), .O(new_n3221));
  nor2 g03028(.a(new_n3019), .b(new_n3012), .O(new_n3222));
  nor2 g03029(.a(new_n3222), .b(new_n3221), .O(new_n3223));
  inv1 g03030(.a(new_n3221), .O(new_n3224));
  inv1 g03031(.a(new_n3222), .O(new_n3225));
  nor2 g03032(.a(new_n3225), .b(new_n3224), .O(new_n3226));
  nor2 g03033(.a(new_n3226), .b(new_n3223), .O(new_n3227));
  inv1 g03034(.a(new_n3227), .O(new_n3228));
  nor2 g03035(.a(new_n2826), .b(new_n196), .O(new_n3229));
  inv1 g03036(.a(new_n3229), .O(new_n3230));
  inv1 g03037(.a(\a[33] ), .O(new_n3231));
  nor2 g03038(.a(new_n3231), .b(new_n198), .O(new_n3232));
  nor2 g03039(.a(new_n1493), .b(new_n502), .O(new_n3233));
  nor2 g03040(.a(new_n3233), .b(new_n3232), .O(new_n3234));
  nor2 g03041(.a(new_n3231), .b(new_n502), .O(new_n3235));
  inv1 g03042(.a(new_n3235), .O(new_n3236));
  nor2 g03043(.a(new_n3236), .b(new_n1504), .O(new_n3237));
  nor2 g03044(.a(new_n3237), .b(new_n3234), .O(new_n3238));
  nor2 g03045(.a(new_n3238), .b(new_n3230), .O(new_n3239));
  inv1 g03046(.a(new_n3238), .O(new_n3240));
  nor2 g03047(.a(new_n3240), .b(new_n3229), .O(new_n3241));
  nor2 g03048(.a(new_n3241), .b(new_n3239), .O(new_n3242));
  nor2 g03049(.a(new_n3242), .b(new_n3228), .O(new_n3243));
  inv1 g03050(.a(new_n3242), .O(new_n3244));
  nor2 g03051(.a(new_n3244), .b(new_n3227), .O(new_n3245));
  nor2 g03052(.a(new_n3245), .b(new_n3243), .O(new_n3246));
  nor2 g03053(.a(new_n3246), .b(new_n3220), .O(new_n3247));
  inv1 g03054(.a(new_n3220), .O(new_n3248));
  inv1 g03055(.a(new_n3246), .O(new_n3249));
  nor2 g03056(.a(new_n3249), .b(new_n3248), .O(new_n3250));
  nor2 g03057(.a(new_n3250), .b(new_n3247), .O(new_n3251));
  inv1 g03058(.a(new_n3251), .O(new_n3252));
  nor2 g03059(.a(new_n941), .b(new_n847), .O(new_n3253));
  nor2 g03060(.a(new_n1086), .b(new_n800), .O(new_n3254));
  nor2 g03061(.a(new_n3254), .b(new_n3253), .O(new_n3255));
  nor2 g03062(.a(new_n1086), .b(new_n847), .O(new_n3256));
  inv1 g03063(.a(new_n3256), .O(new_n3257));
  nor2 g03064(.a(new_n3257), .b(new_n2895), .O(new_n3258));
  nor2 g03065(.a(new_n3258), .b(new_n3255), .O(new_n3259));
  nor2 g03066(.a(new_n3259), .b(new_n2881), .O(new_n3260));
  inv1 g03067(.a(new_n3259), .O(new_n3261));
  nor2 g03068(.a(new_n3261), .b(new_n2880), .O(new_n3262));
  nor2 g03069(.a(new_n3262), .b(new_n3260), .O(new_n3263));
  nor2 g03070(.a(new_n2660), .b(new_n203), .O(new_n3264));
  inv1 g03071(.a(new_n3264), .O(new_n3265));
  nor2 g03072(.a(new_n2506), .b(new_n214), .O(new_n3266));
  nor2 g03073(.a(new_n1736), .b(new_n363), .O(new_n3267));
  nor2 g03074(.a(new_n3267), .b(new_n3266), .O(new_n3268));
  inv1 g03075(.a(new_n3266), .O(new_n3269));
  inv1 g03076(.a(new_n3267), .O(new_n3270));
  nor2 g03077(.a(new_n3270), .b(new_n3269), .O(new_n3271));
  nor2 g03078(.a(new_n3271), .b(new_n3268), .O(new_n3272));
  nor2 g03079(.a(new_n3272), .b(new_n3265), .O(new_n3273));
  inv1 g03080(.a(new_n3272), .O(new_n3274));
  nor2 g03081(.a(new_n3274), .b(new_n3264), .O(new_n3275));
  nor2 g03082(.a(new_n3275), .b(new_n3273), .O(new_n3276));
  nor2 g03083(.a(new_n1903), .b(new_n322), .O(new_n3277));
  nor2 g03084(.a(new_n2184), .b(new_n257), .O(new_n3278));
  nor2 g03085(.a(new_n3278), .b(new_n3277), .O(new_n3279));
  nor2 g03086(.a(new_n2184), .b(new_n322), .O(new_n3280));
  inv1 g03087(.a(new_n3280), .O(new_n3281));
  nor2 g03088(.a(new_n3281), .b(new_n2890), .O(new_n3282));
  nor2 g03089(.a(new_n3282), .b(new_n3279), .O(new_n3283));
  nor2 g03090(.a(new_n3283), .b(new_n3015), .O(new_n3284));
  inv1 g03091(.a(new_n3283), .O(new_n3285));
  nor2 g03092(.a(new_n3285), .b(new_n3014), .O(new_n3286));
  nor2 g03093(.a(new_n3286), .b(new_n3284), .O(new_n3287));
  nor2 g03094(.a(new_n3287), .b(new_n3276), .O(new_n3288));
  inv1 g03095(.a(new_n3276), .O(new_n3289));
  inv1 g03096(.a(new_n3287), .O(new_n3290));
  nor2 g03097(.a(new_n3290), .b(new_n3289), .O(new_n3291));
  nor2 g03098(.a(new_n3291), .b(new_n3288), .O(new_n3292));
  inv1 g03099(.a(new_n3292), .O(new_n3293));
  nor2 g03100(.a(new_n3293), .b(new_n3263), .O(new_n3294));
  inv1 g03101(.a(new_n3263), .O(new_n3295));
  nor2 g03102(.a(new_n3292), .b(new_n3295), .O(new_n3296));
  nor2 g03103(.a(new_n3296), .b(new_n3294), .O(new_n3297));
  inv1 g03104(.a(new_n3297), .O(new_n3298));
  nor2 g03105(.a(new_n3298), .b(new_n3252), .O(new_n3299));
  nor2 g03106(.a(new_n3297), .b(new_n3251), .O(new_n3300));
  nor2 g03107(.a(new_n3300), .b(new_n3299), .O(new_n3301));
  inv1 g03108(.a(new_n3301), .O(new_n3302));
  nor2 g03109(.a(new_n3302), .b(new_n3207), .O(new_n3303));
  nor2 g03110(.a(new_n3301), .b(new_n3206), .O(new_n3304));
  nor2 g03111(.a(new_n3304), .b(new_n3303), .O(new_n3305));
  inv1 g03112(.a(new_n3305), .O(new_n3306));
  nor2 g03113(.a(new_n3137), .b(new_n3132), .O(new_n3307));
  inv1 g03114(.a(new_n3307), .O(new_n3308));
  nor2 g03115(.a(new_n1425), .b(new_n569), .O(new_n3309));
  inv1 g03116(.a(new_n3309), .O(new_n3310));
  nor2 g03117(.a(new_n1199), .b(new_n699), .O(new_n3311));
  nor2 g03118(.a(new_n3311), .b(new_n3074), .O(new_n3312));
  nor2 g03119(.a(new_n1297), .b(new_n699), .O(new_n3313));
  inv1 g03120(.a(new_n3313), .O(new_n3314));
  nor2 g03121(.a(new_n3314), .b(new_n2846), .O(new_n3315));
  nor2 g03122(.a(new_n3315), .b(new_n3312), .O(new_n3316));
  nor2 g03123(.a(new_n3316), .b(new_n3310), .O(new_n3317));
  inv1 g03124(.a(new_n3316), .O(new_n3318));
  nor2 g03125(.a(new_n3318), .b(new_n3309), .O(new_n3319));
  nor2 g03126(.a(new_n3319), .b(new_n3317), .O(new_n3320));
  nor2 g03127(.a(new_n1647), .b(new_n438), .O(new_n3321));
  nor2 g03128(.a(new_n3321), .b(new_n3126), .O(new_n3322));
  inv1 g03129(.a(new_n3126), .O(new_n3323));
  inv1 g03130(.a(new_n3321), .O(new_n3324));
  nor2 g03131(.a(new_n3324), .b(new_n3323), .O(new_n3325));
  nor2 g03132(.a(new_n3325), .b(new_n3322), .O(new_n3326));
  inv1 g03133(.a(new_n3326), .O(new_n3327));
  nor2 g03134(.a(new_n3057), .b(new_n194), .O(new_n3328));
  inv1 g03135(.a(new_n3328), .O(new_n3329));
  nor2 g03136(.a(new_n3329), .b(new_n941), .O(new_n3330));
  nor2 g03137(.a(new_n3328), .b(\a[17] ), .O(new_n3331));
  nor2 g03138(.a(new_n3331), .b(new_n3330), .O(new_n3332));
  inv1 g03139(.a(new_n3332), .O(new_n3333));
  nor2 g03140(.a(new_n3333), .b(new_n3327), .O(new_n3334));
  nor2 g03141(.a(new_n3332), .b(new_n3326), .O(new_n3335));
  nor2 g03142(.a(new_n3335), .b(new_n3334), .O(new_n3336));
  inv1 g03143(.a(new_n3336), .O(new_n3337));
  nor2 g03144(.a(new_n3337), .b(new_n3320), .O(new_n3338));
  inv1 g03145(.a(new_n3320), .O(new_n3339));
  nor2 g03146(.a(new_n3336), .b(new_n3339), .O(new_n3340));
  nor2 g03147(.a(new_n3340), .b(new_n3338), .O(new_n3341));
  nor2 g03148(.a(new_n3341), .b(new_n3308), .O(new_n3342));
  inv1 g03149(.a(new_n3341), .O(new_n3343));
  nor2 g03150(.a(new_n3343), .b(new_n3307), .O(new_n3344));
  nor2 g03151(.a(new_n3344), .b(new_n3342), .O(new_n3345));
  nor2 g03152(.a(new_n3160), .b(new_n3154), .O(new_n3346));
  inv1 g03153(.a(new_n3346), .O(new_n3347));
  nor2 g03154(.a(new_n3347), .b(new_n3345), .O(new_n3348));
  inv1 g03155(.a(new_n3345), .O(new_n3349));
  nor2 g03156(.a(new_n3346), .b(new_n3349), .O(new_n3350));
  nor2 g03157(.a(new_n3350), .b(new_n3348), .O(new_n3351));
  nor2 g03158(.a(new_n3146), .b(new_n3141), .O(new_n3352));
  inv1 g03159(.a(new_n3352), .O(new_n3353));
  nor2 g03160(.a(new_n3353), .b(new_n3351), .O(new_n3354));
  inv1 g03161(.a(new_n3351), .O(new_n3355));
  nor2 g03162(.a(new_n3352), .b(new_n3355), .O(new_n3356));
  nor2 g03163(.a(new_n3356), .b(new_n3354), .O(new_n3357));
  inv1 g03164(.a(new_n3357), .O(new_n3358));
  nor2 g03165(.a(new_n3169), .b(new_n3166), .O(new_n3359));
  nor2 g03166(.a(new_n3359), .b(new_n3358), .O(new_n3360));
  inv1 g03167(.a(new_n3359), .O(new_n3361));
  nor2 g03168(.a(new_n3361), .b(new_n3357), .O(new_n3362));
  nor2 g03169(.a(new_n3362), .b(new_n3360), .O(new_n3363));
  inv1 g03170(.a(new_n3363), .O(new_n3364));
  nor2 g03171(.a(new_n3364), .b(new_n3306), .O(new_n3365));
  nor2 g03172(.a(new_n3363), .b(new_n3305), .O(new_n3366));
  nor2 g03173(.a(new_n3366), .b(new_n3365), .O(new_n3367));
  nor2 g03174(.a(new_n3173), .b(new_n3102), .O(new_n3368));
  inv1 g03175(.a(new_n3368), .O(new_n3369));
  nor2 g03176(.a(new_n3369), .b(new_n3367), .O(new_n3370));
  inv1 g03177(.a(new_n3367), .O(new_n3371));
  nor2 g03178(.a(new_n3368), .b(new_n3371), .O(new_n3372));
  nor2 g03179(.a(new_n3372), .b(new_n3370), .O(new_n3373));
  inv1 g03180(.a(new_n3373), .O(new_n3374));
  nor2 g03181(.a(new_n3183), .b(new_n3179), .O(new_n3375));
  nor2 g03182(.a(new_n3375), .b(new_n3374), .O(new_n3376));
  inv1 g03183(.a(new_n3375), .O(new_n3377));
  nor2 g03184(.a(new_n3377), .b(new_n3373), .O(new_n3378));
  nor2 g03185(.a(new_n3378), .b(new_n3376), .O(new_n3379));
  inv1 g03186(.a(new_n3379), .O(\asquared[34] ));
  nor2 g03187(.a(new_n3365), .b(new_n3360), .O(new_n3381));
  nor2 g03188(.a(new_n3356), .b(new_n3350), .O(new_n3382));
  inv1 g03189(.a(new_n3382), .O(new_n3383));
  nor2 g03190(.a(new_n3275), .b(new_n3268), .O(new_n3384));
  nor2 g03191(.a(new_n3241), .b(new_n3234), .O(new_n3385));
  nor2 g03192(.a(new_n3385), .b(new_n3384), .O(new_n3386));
  inv1 g03193(.a(new_n3384), .O(new_n3387));
  inv1 g03194(.a(new_n3385), .O(new_n3388));
  nor2 g03195(.a(new_n3388), .b(new_n3387), .O(new_n3389));
  nor2 g03196(.a(new_n3389), .b(new_n3386), .O(new_n3390));
  nor2 g03197(.a(new_n3286), .b(new_n3279), .O(new_n3391));
  nor2 g03198(.a(new_n3391), .b(new_n3390), .O(new_n3392));
  inv1 g03199(.a(new_n3390), .O(new_n3393));
  inv1 g03200(.a(new_n3391), .O(new_n3394));
  nor2 g03201(.a(new_n3394), .b(new_n3393), .O(new_n3395));
  nor2 g03202(.a(new_n3395), .b(new_n3392), .O(new_n3396));
  inv1 g03203(.a(new_n3396), .O(new_n3397));
  nor2 g03204(.a(new_n3294), .b(new_n3288), .O(new_n3398));
  inv1 g03205(.a(new_n3330), .O(new_n3399));
  nor2 g03206(.a(new_n3231), .b(new_n194), .O(new_n3400));
  nor2 g03207(.a(new_n3400), .b(new_n3256), .O(new_n3401));
  inv1 g03208(.a(new_n3400), .O(new_n3402));
  nor2 g03209(.a(new_n3402), .b(new_n3257), .O(new_n3403));
  nor2 g03210(.a(new_n3403), .b(new_n3401), .O(new_n3404));
  inv1 g03211(.a(new_n3404), .O(new_n3405));
  nor2 g03212(.a(new_n3405), .b(new_n3399), .O(new_n3406));
  nor2 g03213(.a(new_n3404), .b(new_n3330), .O(new_n3407));
  nor2 g03214(.a(new_n3407), .b(new_n3406), .O(new_n3408));
  inv1 g03215(.a(new_n3408), .O(new_n3409));
  nor2 g03216(.a(new_n3262), .b(new_n3255), .O(new_n3410));
  inv1 g03217(.a(new_n3410), .O(new_n3411));
  nor2 g03218(.a(new_n3411), .b(new_n3409), .O(new_n3412));
  nor2 g03219(.a(new_n3410), .b(new_n3408), .O(new_n3413));
  nor2 g03220(.a(new_n3413), .b(new_n3412), .O(new_n3414));
  inv1 g03221(.a(new_n3414), .O(new_n3415));
  nor2 g03222(.a(new_n3415), .b(new_n3398), .O(new_n3416));
  inv1 g03223(.a(new_n3398), .O(new_n3417));
  nor2 g03224(.a(new_n3414), .b(new_n3417), .O(new_n3418));
  nor2 g03225(.a(new_n3418), .b(new_n3416), .O(new_n3419));
  inv1 g03226(.a(new_n3419), .O(new_n3420));
  nor2 g03227(.a(new_n3420), .b(new_n3397), .O(new_n3421));
  nor2 g03228(.a(new_n3419), .b(new_n3396), .O(new_n3422));
  nor2 g03229(.a(new_n3422), .b(new_n3421), .O(new_n3423));
  inv1 g03230(.a(new_n3423), .O(new_n3424));
  nor2 g03231(.a(new_n3344), .b(new_n3338), .O(new_n3425));
  inv1 g03232(.a(new_n3425), .O(new_n3426));
  nor2 g03233(.a(new_n3334), .b(new_n3325), .O(new_n3427));
  inv1 g03234(.a(new_n3427), .O(new_n3428));
  nor2 g03235(.a(new_n3319), .b(new_n3312), .O(new_n3429));
  nor2 g03236(.a(new_n3429), .b(new_n3428), .O(new_n3430));
  inv1 g03237(.a(new_n3429), .O(new_n3431));
  nor2 g03238(.a(new_n3431), .b(new_n3427), .O(new_n3432));
  nor2 g03239(.a(new_n3432), .b(new_n3430), .O(new_n3433));
  inv1 g03240(.a(new_n3433), .O(new_n3434));
  nor2 g03241(.a(new_n1647), .b(new_n502), .O(new_n3435));
  nor2 g03242(.a(new_n1493), .b(new_n569), .O(new_n3436));
  nor2 g03243(.a(new_n3436), .b(new_n3435), .O(new_n3437));
  inv1 g03244(.a(new_n3233), .O(new_n3438));
  nor2 g03245(.a(new_n1647), .b(new_n569), .O(new_n3439));
  inv1 g03246(.a(new_n3439), .O(new_n3440));
  nor2 g03247(.a(new_n3440), .b(new_n3438), .O(new_n3441));
  nor2 g03248(.a(new_n3441), .b(new_n3437), .O(new_n3442));
  nor2 g03249(.a(new_n3442), .b(new_n3062), .O(new_n3443));
  inv1 g03250(.a(new_n3442), .O(new_n3444));
  nor2 g03251(.a(new_n3444), .b(new_n3061), .O(new_n3445));
  nor2 g03252(.a(new_n3445), .b(new_n3443), .O(new_n3446));
  nor2 g03253(.a(new_n3446), .b(new_n3434), .O(new_n3447));
  inv1 g03254(.a(new_n3446), .O(new_n3448));
  nor2 g03255(.a(new_n3448), .b(new_n3433), .O(new_n3449));
  nor2 g03256(.a(new_n3449), .b(new_n3447), .O(new_n3450));
  nor2 g03257(.a(new_n3450), .b(new_n3426), .O(new_n3451));
  inv1 g03258(.a(new_n3450), .O(new_n3452));
  nor2 g03259(.a(new_n3452), .b(new_n3425), .O(new_n3453));
  nor2 g03260(.a(new_n3453), .b(new_n3451), .O(new_n3454));
  inv1 g03261(.a(new_n3454), .O(new_n3455));
  nor2 g03262(.a(new_n2433), .b(new_n257), .O(new_n3456));
  inv1 g03263(.a(new_n3456), .O(new_n3457));
  nor2 g03264(.a(new_n2184), .b(new_n295), .O(new_n3458));
  nor2 g03265(.a(new_n3458), .b(new_n2577), .O(new_n3459));
  nor2 g03266(.a(new_n3281), .b(new_n2881), .O(new_n3460));
  nor2 g03267(.a(new_n3460), .b(new_n3459), .O(new_n3461));
  nor2 g03268(.a(new_n3461), .b(new_n3457), .O(new_n3462));
  inv1 g03269(.a(new_n3461), .O(new_n3463));
  nor2 g03270(.a(new_n3463), .b(new_n3456), .O(new_n3464));
  nor2 g03271(.a(new_n3464), .b(new_n3462), .O(new_n3465));
  inv1 g03272(.a(new_n3465), .O(new_n3466));
  nor2 g03273(.a(new_n1425), .b(new_n613), .O(new_n3467));
  inv1 g03274(.a(new_n3467), .O(new_n3468));
  nor2 g03275(.a(new_n1199), .b(new_n800), .O(new_n3469));
  nor2 g03276(.a(new_n3469), .b(new_n3313), .O(new_n3470));
  inv1 g03277(.a(new_n3311), .O(new_n3471));
  nor2 g03278(.a(new_n1297), .b(new_n800), .O(new_n3472));
  inv1 g03279(.a(new_n3472), .O(new_n3473));
  nor2 g03280(.a(new_n3473), .b(new_n3471), .O(new_n3474));
  nor2 g03281(.a(new_n3474), .b(new_n3470), .O(new_n3475));
  nor2 g03282(.a(new_n3475), .b(new_n3468), .O(new_n3476));
  inv1 g03283(.a(new_n3475), .O(new_n3477));
  nor2 g03284(.a(new_n3477), .b(new_n3467), .O(new_n3478));
  nor2 g03285(.a(new_n3478), .b(new_n3476), .O(new_n3479));
  nor2 g03286(.a(new_n1736), .b(new_n438), .O(new_n3480));
  inv1 g03287(.a(new_n3480), .O(new_n3481));
  nor2 g03288(.a(new_n2506), .b(new_n229), .O(new_n3482));
  nor2 g03289(.a(new_n1903), .b(new_n363), .O(new_n3483));
  nor2 g03290(.a(new_n3483), .b(new_n3482), .O(new_n3484));
  inv1 g03291(.a(new_n3482), .O(new_n3485));
  inv1 g03292(.a(new_n3483), .O(new_n3486));
  nor2 g03293(.a(new_n3486), .b(new_n3485), .O(new_n3487));
  nor2 g03294(.a(new_n3487), .b(new_n3484), .O(new_n3488));
  nor2 g03295(.a(new_n3488), .b(new_n3481), .O(new_n3489));
  inv1 g03296(.a(new_n3488), .O(new_n3490));
  nor2 g03297(.a(new_n3490), .b(new_n3480), .O(new_n3491));
  nor2 g03298(.a(new_n3491), .b(new_n3489), .O(new_n3492));
  nor2 g03299(.a(new_n3492), .b(new_n3479), .O(new_n3493));
  inv1 g03300(.a(new_n3479), .O(new_n3494));
  inv1 g03301(.a(new_n3492), .O(new_n3495));
  nor2 g03302(.a(new_n3495), .b(new_n3494), .O(new_n3496));
  nor2 g03303(.a(new_n3496), .b(new_n3493), .O(new_n3497));
  nor2 g03304(.a(new_n3497), .b(new_n3466), .O(new_n3498));
  inv1 g03305(.a(new_n3497), .O(new_n3499));
  nor2 g03306(.a(new_n3499), .b(new_n3465), .O(new_n3500));
  nor2 g03307(.a(new_n3500), .b(new_n3498), .O(new_n3501));
  inv1 g03308(.a(new_n3501), .O(new_n3502));
  nor2 g03309(.a(new_n3502), .b(new_n3455), .O(new_n3503));
  nor2 g03310(.a(new_n3501), .b(new_n3454), .O(new_n3504));
  nor2 g03311(.a(new_n3504), .b(new_n3503), .O(new_n3505));
  inv1 g03312(.a(new_n3505), .O(new_n3506));
  nor2 g03313(.a(new_n3506), .b(new_n3424), .O(new_n3507));
  nor2 g03314(.a(new_n3505), .b(new_n3423), .O(new_n3508));
  nor2 g03315(.a(new_n3508), .b(new_n3507), .O(new_n3509));
  nor2 g03316(.a(new_n3509), .b(new_n3383), .O(new_n3510));
  inv1 g03317(.a(new_n3509), .O(new_n3511));
  nor2 g03318(.a(new_n3511), .b(new_n3382), .O(new_n3512));
  nor2 g03319(.a(new_n3512), .b(new_n3510), .O(new_n3513));
  inv1 g03320(.a(new_n3513), .O(new_n3514));
  nor2 g03321(.a(new_n3303), .b(new_n3203), .O(new_n3515));
  inv1 g03322(.a(new_n3515), .O(new_n3516));
  nor2 g03323(.a(new_n3299), .b(new_n3250), .O(new_n3517));
  inv1 g03324(.a(new_n3517), .O(new_n3518));
  nor2 g03325(.a(new_n3199), .b(new_n3193), .O(new_n3519));
  inv1 g03326(.a(new_n3519), .O(new_n3520));
  nor2 g03327(.a(new_n3520), .b(new_n3518), .O(new_n3521));
  nor2 g03328(.a(new_n3519), .b(new_n3517), .O(new_n3522));
  nor2 g03329(.a(new_n3522), .b(new_n3521), .O(new_n3523));
  inv1 g03330(.a(new_n3523), .O(new_n3524));
  nor2 g03331(.a(new_n3219), .b(new_n3213), .O(new_n3525));
  nor2 g03332(.a(new_n2826), .b(new_n203), .O(new_n3526));
  nor2 g03333(.a(new_n2660), .b(new_n214), .O(new_n3527));
  nor2 g03334(.a(new_n3527), .b(new_n3526), .O(new_n3528));
  nor2 g03335(.a(new_n2826), .b(new_n214), .O(new_n3529));
  inv1 g03336(.a(new_n3529), .O(new_n3530));
  nor2 g03337(.a(new_n3530), .b(new_n3265), .O(new_n3531));
  nor2 g03338(.a(new_n3531), .b(new_n3528), .O(new_n3532));
  inv1 g03339(.a(\a[34] ), .O(new_n3533));
  nor2 g03340(.a(new_n3533), .b(new_n198), .O(new_n3534));
  inv1 g03341(.a(new_n3534), .O(new_n3535));
  nor2 g03342(.a(new_n3535), .b(new_n3532), .O(new_n3536));
  inv1 g03343(.a(new_n3532), .O(new_n3537));
  nor2 g03344(.a(new_n3534), .b(new_n3537), .O(new_n3538));
  nor2 g03345(.a(new_n3538), .b(new_n3536), .O(new_n3539));
  nor2 g03346(.a(new_n3539), .b(new_n3525), .O(new_n3540));
  inv1 g03347(.a(new_n3525), .O(new_n3541));
  inv1 g03348(.a(new_n3539), .O(new_n3542));
  nor2 g03349(.a(new_n3542), .b(new_n3541), .O(new_n3543));
  nor2 g03350(.a(new_n3543), .b(new_n3540), .O(new_n3544));
  inv1 g03351(.a(new_n3544), .O(new_n3545));
  nor2 g03352(.a(new_n3243), .b(new_n3226), .O(new_n3546));
  nor2 g03353(.a(new_n3546), .b(new_n3545), .O(new_n3547));
  inv1 g03354(.a(new_n3546), .O(new_n3548));
  nor2 g03355(.a(new_n3548), .b(new_n3544), .O(new_n3549));
  nor2 g03356(.a(new_n3549), .b(new_n3547), .O(new_n3550));
  inv1 g03357(.a(new_n3550), .O(new_n3551));
  nor2 g03358(.a(new_n3551), .b(new_n3524), .O(new_n3552));
  nor2 g03359(.a(new_n3550), .b(new_n3523), .O(new_n3553));
  nor2 g03360(.a(new_n3553), .b(new_n3552), .O(new_n3554));
  nor2 g03361(.a(new_n3554), .b(new_n3516), .O(new_n3555));
  inv1 g03362(.a(new_n3554), .O(new_n3556));
  nor2 g03363(.a(new_n3556), .b(new_n3515), .O(new_n3557));
  nor2 g03364(.a(new_n3557), .b(new_n3555), .O(new_n3558));
  inv1 g03365(.a(new_n3558), .O(new_n3559));
  nor2 g03366(.a(new_n3559), .b(new_n3514), .O(new_n3560));
  nor2 g03367(.a(new_n3558), .b(new_n3513), .O(new_n3561));
  nor2 g03368(.a(new_n3561), .b(new_n3560), .O(new_n3562));
  inv1 g03369(.a(new_n3562), .O(new_n3563));
  nor2 g03370(.a(new_n3563), .b(new_n3381), .O(new_n3564));
  inv1 g03371(.a(new_n3381), .O(new_n3565));
  nor2 g03372(.a(new_n3562), .b(new_n3565), .O(new_n3566));
  nor2 g03373(.a(new_n3566), .b(new_n3564), .O(new_n3567));
  inv1 g03374(.a(new_n3567), .O(new_n3568));
  nor2 g03375(.a(new_n3376), .b(new_n3370), .O(new_n3569));
  nor2 g03376(.a(new_n3569), .b(new_n3568), .O(new_n3570));
  inv1 g03377(.a(new_n3569), .O(new_n3571));
  nor2 g03378(.a(new_n3571), .b(new_n3567), .O(new_n3572));
  nor2 g03379(.a(new_n3572), .b(new_n3570), .O(new_n3573));
  inv1 g03380(.a(new_n3573), .O(\asquared[35] ));
  nor2 g03381(.a(new_n3560), .b(new_n3557), .O(new_n3575));
  inv1 g03382(.a(new_n3575), .O(new_n3576));
  nor2 g03383(.a(new_n3512), .b(new_n3507), .O(new_n3577));
  inv1 g03384(.a(new_n3577), .O(new_n3578));
  nor2 g03385(.a(new_n3395), .b(new_n3389), .O(new_n3579));
  inv1 g03386(.a(new_n3579), .O(new_n3580));
  nor2 g03387(.a(new_n3412), .b(new_n3406), .O(new_n3581));
  inv1 g03388(.a(new_n3581), .O(new_n3582));
  nor2 g03389(.a(new_n3582), .b(new_n3580), .O(new_n3583));
  nor2 g03390(.a(new_n3581), .b(new_n3579), .O(new_n3584));
  nor2 g03391(.a(new_n3584), .b(new_n3583), .O(new_n3585));
  nor2 g03392(.a(new_n3447), .b(new_n3432), .O(new_n3586));
  inv1 g03393(.a(new_n3586), .O(new_n3587));
  nor2 g03394(.a(new_n3587), .b(new_n3585), .O(new_n3588));
  inv1 g03395(.a(new_n3585), .O(new_n3589));
  nor2 g03396(.a(new_n3586), .b(new_n3589), .O(new_n3590));
  nor2 g03397(.a(new_n3590), .b(new_n3588), .O(new_n3591));
  nor2 g03398(.a(new_n3421), .b(new_n3416), .O(new_n3592));
  inv1 g03399(.a(new_n3592), .O(new_n3593));
  nor2 g03400(.a(new_n3593), .b(new_n3591), .O(new_n3594));
  inv1 g03401(.a(new_n3591), .O(new_n3595));
  nor2 g03402(.a(new_n3592), .b(new_n3595), .O(new_n3596));
  nor2 g03403(.a(new_n3596), .b(new_n3594), .O(new_n3597));
  inv1 g03404(.a(new_n3597), .O(new_n3598));
  nor2 g03405(.a(new_n3503), .b(new_n3453), .O(new_n3599));
  nor2 g03406(.a(new_n3599), .b(new_n3598), .O(new_n3600));
  inv1 g03407(.a(new_n3599), .O(new_n3601));
  nor2 g03408(.a(new_n3601), .b(new_n3597), .O(new_n3602));
  nor2 g03409(.a(new_n3602), .b(new_n3600), .O(new_n3603));
  nor2 g03410(.a(new_n3603), .b(new_n3578), .O(new_n3604));
  inv1 g03411(.a(new_n3603), .O(new_n3605));
  nor2 g03412(.a(new_n3605), .b(new_n3577), .O(new_n3606));
  nor2 g03413(.a(new_n3606), .b(new_n3604), .O(new_n3607));
  nor2 g03414(.a(new_n3552), .b(new_n3522), .O(new_n3608));
  nor2 g03415(.a(new_n3445), .b(new_n3437), .O(new_n3609));
  nor2 g03416(.a(new_n3478), .b(new_n3470), .O(new_n3610));
  nor2 g03417(.a(new_n3610), .b(new_n3609), .O(new_n3611));
  inv1 g03418(.a(new_n3609), .O(new_n3612));
  inv1 g03419(.a(new_n3610), .O(new_n3613));
  nor2 g03420(.a(new_n3613), .b(new_n3612), .O(new_n3614));
  nor2 g03421(.a(new_n3614), .b(new_n3611), .O(new_n3615));
  nor2 g03422(.a(new_n3538), .b(new_n3528), .O(new_n3616));
  nor2 g03423(.a(new_n3616), .b(new_n3615), .O(new_n3617));
  inv1 g03424(.a(new_n3615), .O(new_n3618));
  inv1 g03425(.a(new_n3616), .O(new_n3619));
  nor2 g03426(.a(new_n3619), .b(new_n3618), .O(new_n3620));
  nor2 g03427(.a(new_n3620), .b(new_n3617), .O(new_n3621));
  inv1 g03428(.a(new_n3621), .O(new_n3622));
  nor2 g03429(.a(new_n1131), .b(new_n3533), .O(new_n3623));
  nor2 g03430(.a(new_n3533), .b(new_n194), .O(new_n3624));
  nor2 g03431(.a(new_n3624), .b(\a[18] ), .O(new_n3625));
  nor2 g03432(.a(new_n3625), .b(new_n3623), .O(new_n3626));
  nor2 g03433(.a(new_n3464), .b(new_n3459), .O(new_n3627));
  nor2 g03434(.a(new_n3627), .b(new_n3626), .O(new_n3628));
  inv1 g03435(.a(new_n3626), .O(new_n3629));
  inv1 g03436(.a(new_n3627), .O(new_n3630));
  nor2 g03437(.a(new_n3630), .b(new_n3629), .O(new_n3631));
  nor2 g03438(.a(new_n3631), .b(new_n3628), .O(new_n3632));
  inv1 g03439(.a(new_n3632), .O(new_n3633));
  nor2 g03440(.a(new_n3491), .b(new_n3484), .O(new_n3634));
  inv1 g03441(.a(new_n3634), .O(new_n3635));
  nor2 g03442(.a(new_n3635), .b(new_n3633), .O(new_n3636));
  nor2 g03443(.a(new_n3634), .b(new_n3632), .O(new_n3637));
  nor2 g03444(.a(new_n3637), .b(new_n3636), .O(new_n3638));
  inv1 g03445(.a(new_n3638), .O(new_n3639));
  nor2 g03446(.a(new_n3500), .b(new_n3493), .O(new_n3640));
  nor2 g03447(.a(new_n3640), .b(new_n3639), .O(new_n3641));
  inv1 g03448(.a(new_n3640), .O(new_n3642));
  nor2 g03449(.a(new_n3642), .b(new_n3638), .O(new_n3643));
  nor2 g03450(.a(new_n3643), .b(new_n3641), .O(new_n3644));
  inv1 g03451(.a(new_n3644), .O(new_n3645));
  nor2 g03452(.a(new_n3645), .b(new_n3622), .O(new_n3646));
  nor2 g03453(.a(new_n3644), .b(new_n3621), .O(new_n3647));
  nor2 g03454(.a(new_n3647), .b(new_n3646), .O(new_n3648));
  inv1 g03455(.a(new_n3648), .O(new_n3649));
  nor2 g03456(.a(new_n3649), .b(new_n3608), .O(new_n3650));
  inv1 g03457(.a(new_n3608), .O(new_n3651));
  nor2 g03458(.a(new_n3648), .b(new_n3651), .O(new_n3652));
  nor2 g03459(.a(new_n3652), .b(new_n3650), .O(new_n3653));
  inv1 g03460(.a(new_n3653), .O(new_n3654));
  nor2 g03461(.a(new_n3547), .b(new_n3540), .O(new_n3655));
  inv1 g03462(.a(new_n3655), .O(new_n3656));
  nor2 g03463(.a(new_n2121), .b(new_n363), .O(new_n3657));
  nor2 g03464(.a(new_n1903), .b(new_n438), .O(new_n3658));
  nor2 g03465(.a(new_n3658), .b(new_n3657), .O(new_n3659));
  nor2 g03466(.a(new_n2121), .b(new_n438), .O(new_n3660));
  inv1 g03467(.a(new_n3660), .O(new_n3661));
  nor2 g03468(.a(new_n3661), .b(new_n3486), .O(new_n3662));
  nor2 g03469(.a(new_n3662), .b(new_n3659), .O(new_n3663));
  nor2 g03470(.a(new_n3663), .b(new_n3530), .O(new_n3664));
  inv1 g03471(.a(new_n3663), .O(new_n3665));
  nor2 g03472(.a(new_n3665), .b(new_n3529), .O(new_n3666));
  nor2 g03473(.a(new_n3666), .b(new_n3664), .O(new_n3667));
  inv1 g03474(.a(new_n3667), .O(new_n3668));
  nor2 g03475(.a(new_n2660), .b(new_n229), .O(new_n3669));
  nor2 g03476(.a(new_n2506), .b(new_n257), .O(new_n3670));
  nor2 g03477(.a(new_n3670), .b(new_n3280), .O(new_n3671));
  inv1 g03478(.a(new_n3278), .O(new_n3672));
  nor2 g03479(.a(new_n2506), .b(new_n322), .O(new_n3673));
  inv1 g03480(.a(new_n3673), .O(new_n3674));
  nor2 g03481(.a(new_n3674), .b(new_n3672), .O(new_n3675));
  nor2 g03482(.a(new_n3675), .b(new_n3671), .O(new_n3676));
  inv1 g03483(.a(new_n3676), .O(new_n3677));
  nor2 g03484(.a(new_n3677), .b(new_n3669), .O(new_n3678));
  inv1 g03485(.a(new_n3669), .O(new_n3679));
  nor2 g03486(.a(new_n3676), .b(new_n3679), .O(new_n3680));
  nor2 g03487(.a(new_n3680), .b(new_n3678), .O(new_n3681));
  nor2 g03488(.a(new_n2433), .b(new_n295), .O(new_n3682));
  inv1 g03489(.a(new_n3682), .O(new_n3683));
  nor2 g03490(.a(new_n1086), .b(new_n941), .O(new_n3684));
  nor2 g03491(.a(new_n1199), .b(new_n847), .O(new_n3685));
  nor2 g03492(.a(new_n3685), .b(new_n3684), .O(new_n3686));
  inv1 g03493(.a(new_n3684), .O(new_n3687));
  inv1 g03494(.a(new_n3685), .O(new_n3688));
  nor2 g03495(.a(new_n3688), .b(new_n3687), .O(new_n3689));
  nor2 g03496(.a(new_n3689), .b(new_n3686), .O(new_n3690));
  nor2 g03497(.a(new_n3690), .b(new_n3683), .O(new_n3691));
  inv1 g03498(.a(new_n3690), .O(new_n3692));
  nor2 g03499(.a(new_n3692), .b(new_n3682), .O(new_n3693));
  nor2 g03500(.a(new_n3693), .b(new_n3691), .O(new_n3694));
  nor2 g03501(.a(new_n3694), .b(new_n3681), .O(new_n3695));
  inv1 g03502(.a(new_n3681), .O(new_n3696));
  inv1 g03503(.a(new_n3694), .O(new_n3697));
  nor2 g03504(.a(new_n3697), .b(new_n3696), .O(new_n3698));
  nor2 g03505(.a(new_n3698), .b(new_n3695), .O(new_n3699));
  nor2 g03506(.a(new_n3699), .b(new_n3668), .O(new_n3700));
  inv1 g03507(.a(new_n3699), .O(new_n3701));
  nor2 g03508(.a(new_n3701), .b(new_n3667), .O(new_n3702));
  nor2 g03509(.a(new_n3702), .b(new_n3700), .O(new_n3703));
  nor2 g03510(.a(new_n3703), .b(new_n3656), .O(new_n3704));
  inv1 g03511(.a(new_n3703), .O(new_n3705));
  nor2 g03512(.a(new_n3705), .b(new_n3655), .O(new_n3706));
  nor2 g03513(.a(new_n3706), .b(new_n3704), .O(new_n3707));
  inv1 g03514(.a(new_n3707), .O(new_n3708));
  nor2 g03515(.a(new_n1493), .b(new_n613), .O(new_n3709));
  inv1 g03516(.a(new_n3709), .O(new_n3710));
  nor2 g03517(.a(new_n1425), .b(new_n699), .O(new_n3711));
  nor2 g03518(.a(new_n3711), .b(new_n3472), .O(new_n3712));
  nor2 g03519(.a(new_n1425), .b(new_n800), .O(new_n3713));
  inv1 g03520(.a(new_n3713), .O(new_n3714));
  nor2 g03521(.a(new_n3714), .b(new_n3314), .O(new_n3715));
  nor2 g03522(.a(new_n3715), .b(new_n3712), .O(new_n3716));
  nor2 g03523(.a(new_n3716), .b(new_n3710), .O(new_n3717));
  inv1 g03524(.a(new_n3716), .O(new_n3718));
  nor2 g03525(.a(new_n3718), .b(new_n3709), .O(new_n3719));
  nor2 g03526(.a(new_n3719), .b(new_n3717), .O(new_n3720));
  inv1 g03527(.a(new_n3720), .O(new_n3721));
  inv1 g03528(.a(\a[35] ), .O(new_n3722));
  nor2 g03529(.a(new_n3722), .b(new_n198), .O(new_n3723));
  nor2 g03530(.a(new_n3231), .b(new_n196), .O(new_n3724));
  nor2 g03531(.a(new_n3724), .b(new_n3723), .O(new_n3725));
  inv1 g03532(.a(new_n3232), .O(new_n3726));
  nor2 g03533(.a(new_n3722), .b(new_n196), .O(new_n3727));
  inv1 g03534(.a(new_n3727), .O(new_n3728));
  nor2 g03535(.a(new_n3728), .b(new_n3726), .O(new_n3729));
  nor2 g03536(.a(new_n3729), .b(new_n3725), .O(new_n3730));
  inv1 g03537(.a(new_n3730), .O(new_n3731));
  nor2 g03538(.a(new_n3731), .b(new_n3403), .O(new_n3732));
  inv1 g03539(.a(new_n3403), .O(new_n3733));
  nor2 g03540(.a(new_n3730), .b(new_n3733), .O(new_n3734));
  nor2 g03541(.a(new_n3734), .b(new_n3732), .O(new_n3735));
  nor2 g03542(.a(new_n3057), .b(new_n203), .O(new_n3736));
  inv1 g03543(.a(new_n3736), .O(new_n3737));
  nor2 g03544(.a(new_n1736), .b(new_n502), .O(new_n3738));
  nor2 g03545(.a(new_n3738), .b(new_n3439), .O(new_n3739));
  inv1 g03546(.a(new_n3435), .O(new_n3740));
  nor2 g03547(.a(new_n1736), .b(new_n569), .O(new_n3741));
  inv1 g03548(.a(new_n3741), .O(new_n3742));
  nor2 g03549(.a(new_n3742), .b(new_n3740), .O(new_n3743));
  nor2 g03550(.a(new_n3743), .b(new_n3739), .O(new_n3744));
  nor2 g03551(.a(new_n3744), .b(new_n3737), .O(new_n3745));
  inv1 g03552(.a(new_n3744), .O(new_n3746));
  nor2 g03553(.a(new_n3746), .b(new_n3736), .O(new_n3747));
  nor2 g03554(.a(new_n3747), .b(new_n3745), .O(new_n3748));
  nor2 g03555(.a(new_n3748), .b(new_n3735), .O(new_n3749));
  inv1 g03556(.a(new_n3735), .O(new_n3750));
  inv1 g03557(.a(new_n3748), .O(new_n3751));
  nor2 g03558(.a(new_n3751), .b(new_n3750), .O(new_n3752));
  nor2 g03559(.a(new_n3752), .b(new_n3749), .O(new_n3753));
  nor2 g03560(.a(new_n3753), .b(new_n3721), .O(new_n3754));
  inv1 g03561(.a(new_n3753), .O(new_n3755));
  nor2 g03562(.a(new_n3755), .b(new_n3720), .O(new_n3756));
  nor2 g03563(.a(new_n3756), .b(new_n3754), .O(new_n3757));
  inv1 g03564(.a(new_n3757), .O(new_n3758));
  nor2 g03565(.a(new_n3758), .b(new_n3708), .O(new_n3759));
  nor2 g03566(.a(new_n3757), .b(new_n3707), .O(new_n3760));
  nor2 g03567(.a(new_n3760), .b(new_n3759), .O(new_n3761));
  inv1 g03568(.a(new_n3761), .O(new_n3762));
  nor2 g03569(.a(new_n3762), .b(new_n3654), .O(new_n3763));
  nor2 g03570(.a(new_n3761), .b(new_n3653), .O(new_n3764));
  nor2 g03571(.a(new_n3764), .b(new_n3763), .O(new_n3765));
  nor2 g03572(.a(new_n3765), .b(new_n3607), .O(new_n3766));
  inv1 g03573(.a(new_n3607), .O(new_n3767));
  inv1 g03574(.a(new_n3765), .O(new_n3768));
  nor2 g03575(.a(new_n3768), .b(new_n3767), .O(new_n3769));
  nor2 g03576(.a(new_n3769), .b(new_n3766), .O(new_n3770));
  nor2 g03577(.a(new_n3770), .b(new_n3576), .O(new_n3771));
  inv1 g03578(.a(new_n3770), .O(new_n3772));
  nor2 g03579(.a(new_n3772), .b(new_n3575), .O(new_n3773));
  nor2 g03580(.a(new_n3773), .b(new_n3771), .O(new_n3774));
  inv1 g03581(.a(new_n3774), .O(new_n3775));
  nor2 g03582(.a(new_n3570), .b(new_n3566), .O(new_n3776));
  nor2 g03583(.a(new_n3776), .b(new_n3775), .O(new_n3777));
  inv1 g03584(.a(new_n3776), .O(new_n3778));
  nor2 g03585(.a(new_n3778), .b(new_n3774), .O(new_n3779));
  nor2 g03586(.a(new_n3779), .b(new_n3777), .O(new_n3780));
  inv1 g03587(.a(new_n3780), .O(\asquared[36] ));
  nor2 g03588(.a(new_n3769), .b(new_n3606), .O(new_n3782));
  inv1 g03589(.a(new_n3782), .O(new_n3783));
  nor2 g03590(.a(new_n3763), .b(new_n3650), .O(new_n3784));
  nor2 g03591(.a(new_n3620), .b(new_n3614), .O(new_n3785));
  inv1 g03592(.a(new_n3785), .O(new_n3786));
  nor2 g03593(.a(new_n3636), .b(new_n3631), .O(new_n3787));
  inv1 g03594(.a(new_n3787), .O(new_n3788));
  nor2 g03595(.a(new_n3788), .b(new_n3786), .O(new_n3789));
  nor2 g03596(.a(new_n3787), .b(new_n3785), .O(new_n3790));
  nor2 g03597(.a(new_n3790), .b(new_n3789), .O(new_n3791));
  nor2 g03598(.a(new_n3756), .b(new_n3749), .O(new_n3792));
  inv1 g03599(.a(new_n3792), .O(new_n3793));
  nor2 g03600(.a(new_n3793), .b(new_n3791), .O(new_n3794));
  inv1 g03601(.a(new_n3791), .O(new_n3795));
  nor2 g03602(.a(new_n3792), .b(new_n3795), .O(new_n3796));
  nor2 g03603(.a(new_n3796), .b(new_n3794), .O(new_n3797));
  nor2 g03604(.a(new_n3646), .b(new_n3641), .O(new_n3798));
  inv1 g03605(.a(new_n3798), .O(new_n3799));
  nor2 g03606(.a(new_n3799), .b(new_n3797), .O(new_n3800));
  inv1 g03607(.a(new_n3797), .O(new_n3801));
  nor2 g03608(.a(new_n3798), .b(new_n3801), .O(new_n3802));
  nor2 g03609(.a(new_n3802), .b(new_n3800), .O(new_n3803));
  inv1 g03610(.a(new_n3803), .O(new_n3804));
  nor2 g03611(.a(new_n3759), .b(new_n3706), .O(new_n3805));
  nor2 g03612(.a(new_n3805), .b(new_n3804), .O(new_n3806));
  inv1 g03613(.a(new_n3805), .O(new_n3807));
  nor2 g03614(.a(new_n3807), .b(new_n3803), .O(new_n3808));
  nor2 g03615(.a(new_n3808), .b(new_n3806), .O(new_n3809));
  inv1 g03616(.a(new_n3809), .O(new_n3810));
  nor2 g03617(.a(new_n3810), .b(new_n3784), .O(new_n3811));
  inv1 g03618(.a(new_n3784), .O(new_n3812));
  nor2 g03619(.a(new_n3809), .b(new_n3812), .O(new_n3813));
  nor2 g03620(.a(new_n3813), .b(new_n3811), .O(new_n3814));
  inv1 g03621(.a(new_n3814), .O(new_n3815));
  nor2 g03622(.a(new_n3600), .b(new_n3596), .O(new_n3816));
  nor2 g03623(.a(new_n3666), .b(new_n3659), .O(new_n3817));
  nor2 g03624(.a(new_n3678), .b(new_n3671), .O(new_n3818));
  nor2 g03625(.a(new_n3818), .b(new_n3817), .O(new_n3819));
  inv1 g03626(.a(new_n3817), .O(new_n3820));
  inv1 g03627(.a(new_n3818), .O(new_n3821));
  nor2 g03628(.a(new_n3821), .b(new_n3820), .O(new_n3822));
  nor2 g03629(.a(new_n3822), .b(new_n3819), .O(new_n3823));
  nor2 g03630(.a(new_n3693), .b(new_n3686), .O(new_n3824));
  nor2 g03631(.a(new_n3824), .b(new_n3823), .O(new_n3825));
  inv1 g03632(.a(new_n3823), .O(new_n3826));
  inv1 g03633(.a(new_n3824), .O(new_n3827));
  nor2 g03634(.a(new_n3827), .b(new_n3826), .O(new_n3828));
  nor2 g03635(.a(new_n3828), .b(new_n3825), .O(new_n3829));
  inv1 g03636(.a(new_n3829), .O(new_n3830));
  nor2 g03637(.a(new_n3747), .b(new_n3739), .O(new_n3831));
  nor2 g03638(.a(new_n3719), .b(new_n3712), .O(new_n3832));
  nor2 g03639(.a(new_n3832), .b(new_n3831), .O(new_n3833));
  inv1 g03640(.a(new_n3831), .O(new_n3834));
  inv1 g03641(.a(new_n3832), .O(new_n3835));
  nor2 g03642(.a(new_n3835), .b(new_n3834), .O(new_n3836));
  nor2 g03643(.a(new_n3836), .b(new_n3833), .O(new_n3837));
  nor2 g03644(.a(new_n3732), .b(new_n3725), .O(new_n3838));
  nor2 g03645(.a(new_n3838), .b(new_n3837), .O(new_n3839));
  inv1 g03646(.a(new_n3837), .O(new_n3840));
  inv1 g03647(.a(new_n3838), .O(new_n3841));
  nor2 g03648(.a(new_n3841), .b(new_n3840), .O(new_n3842));
  nor2 g03649(.a(new_n3842), .b(new_n3839), .O(new_n3843));
  nor2 g03650(.a(new_n3702), .b(new_n3695), .O(new_n3844));
  inv1 g03651(.a(new_n3844), .O(new_n3845));
  nor2 g03652(.a(new_n3845), .b(new_n3843), .O(new_n3846));
  inv1 g03653(.a(new_n3843), .O(new_n3847));
  nor2 g03654(.a(new_n3844), .b(new_n3847), .O(new_n3848));
  nor2 g03655(.a(new_n3848), .b(new_n3846), .O(new_n3849));
  inv1 g03656(.a(new_n3849), .O(new_n3850));
  nor2 g03657(.a(new_n3850), .b(new_n3830), .O(new_n3851));
  nor2 g03658(.a(new_n3849), .b(new_n3829), .O(new_n3852));
  nor2 g03659(.a(new_n3852), .b(new_n3851), .O(new_n3853));
  inv1 g03660(.a(new_n3853), .O(new_n3854));
  nor2 g03661(.a(new_n3854), .b(new_n3816), .O(new_n3855));
  inv1 g03662(.a(new_n3816), .O(new_n3856));
  nor2 g03663(.a(new_n3853), .b(new_n3856), .O(new_n3857));
  nor2 g03664(.a(new_n3857), .b(new_n3855), .O(new_n3858));
  inv1 g03665(.a(new_n3858), .O(new_n3859));
  nor2 g03666(.a(new_n3590), .b(new_n3584), .O(new_n3860));
  nor2 g03667(.a(new_n1199), .b(new_n941), .O(new_n3861));
  nor2 g03668(.a(new_n3722), .b(new_n194), .O(new_n3862));
  nor2 g03669(.a(new_n3862), .b(new_n3861), .O(new_n3863));
  inv1 g03670(.a(new_n3861), .O(new_n3864));
  inv1 g03671(.a(new_n3862), .O(new_n3865));
  nor2 g03672(.a(new_n3865), .b(new_n3864), .O(new_n3866));
  nor2 g03673(.a(new_n3866), .b(new_n3863), .O(new_n3867));
  inv1 g03674(.a(new_n3867), .O(new_n3868));
  inv1 g03675(.a(new_n3623), .O(new_n3869));
  inv1 g03676(.a(\a[36] ), .O(new_n3870));
  nor2 g03677(.a(new_n3870), .b(new_n198), .O(new_n3871));
  inv1 g03678(.a(new_n3871), .O(new_n3872));
  nor2 g03679(.a(new_n3872), .b(new_n3869), .O(new_n3873));
  nor2 g03680(.a(new_n3871), .b(new_n3623), .O(new_n3874));
  nor2 g03681(.a(new_n3874), .b(new_n3873), .O(new_n3875));
  inv1 g03682(.a(new_n3875), .O(new_n3876));
  nor2 g03683(.a(new_n3876), .b(new_n3868), .O(new_n3877));
  nor2 g03684(.a(new_n3875), .b(new_n3867), .O(new_n3878));
  nor2 g03685(.a(new_n3878), .b(new_n3877), .O(new_n3879));
  inv1 g03686(.a(new_n3879), .O(new_n3880));
  nor2 g03687(.a(new_n1493), .b(new_n699), .O(new_n3881));
  inv1 g03688(.a(new_n3881), .O(new_n3882));
  nor2 g03689(.a(new_n1297), .b(new_n847), .O(new_n3883));
  nor2 g03690(.a(new_n3883), .b(new_n3713), .O(new_n3884));
  nor2 g03691(.a(new_n1425), .b(new_n847), .O(new_n3885));
  inv1 g03692(.a(new_n3885), .O(new_n3886));
  nor2 g03693(.a(new_n3886), .b(new_n3473), .O(new_n3887));
  nor2 g03694(.a(new_n3887), .b(new_n3884), .O(new_n3888));
  nor2 g03695(.a(new_n3888), .b(new_n3882), .O(new_n3889));
  inv1 g03696(.a(new_n3888), .O(new_n3890));
  nor2 g03697(.a(new_n3890), .b(new_n3881), .O(new_n3891));
  nor2 g03698(.a(new_n3891), .b(new_n3889), .O(new_n3892));
  nor2 g03699(.a(new_n3231), .b(new_n203), .O(new_n3893));
  inv1 g03700(.a(new_n3893), .O(new_n3894));
  nor2 g03701(.a(new_n1903), .b(new_n502), .O(new_n3895));
  nor2 g03702(.a(new_n3057), .b(new_n214), .O(new_n3896));
  nor2 g03703(.a(new_n3896), .b(new_n3895), .O(new_n3897));
  inv1 g03704(.a(new_n3895), .O(new_n3898));
  inv1 g03705(.a(new_n3896), .O(new_n3899));
  nor2 g03706(.a(new_n3899), .b(new_n3898), .O(new_n3900));
  nor2 g03707(.a(new_n3900), .b(new_n3897), .O(new_n3901));
  nor2 g03708(.a(new_n3901), .b(new_n3894), .O(new_n3902));
  inv1 g03709(.a(new_n3901), .O(new_n3903));
  nor2 g03710(.a(new_n3903), .b(new_n3893), .O(new_n3904));
  nor2 g03711(.a(new_n3904), .b(new_n3902), .O(new_n3905));
  nor2 g03712(.a(new_n3905), .b(new_n3892), .O(new_n3906));
  inv1 g03713(.a(new_n3892), .O(new_n3907));
  inv1 g03714(.a(new_n3905), .O(new_n3908));
  nor2 g03715(.a(new_n3908), .b(new_n3907), .O(new_n3909));
  nor2 g03716(.a(new_n3909), .b(new_n3906), .O(new_n3910));
  inv1 g03717(.a(new_n3910), .O(new_n3911));
  nor2 g03718(.a(new_n3911), .b(new_n3880), .O(new_n3912));
  nor2 g03719(.a(new_n3910), .b(new_n3879), .O(new_n3913));
  nor2 g03720(.a(new_n3913), .b(new_n3912), .O(new_n3914));
  inv1 g03721(.a(new_n3914), .O(new_n3915));
  nor2 g03722(.a(new_n3915), .b(new_n3860), .O(new_n3916));
  inv1 g03723(.a(new_n3860), .O(new_n3917));
  nor2 g03724(.a(new_n3914), .b(new_n3917), .O(new_n3918));
  nor2 g03725(.a(new_n3918), .b(new_n3916), .O(new_n3919));
  inv1 g03726(.a(new_n3919), .O(new_n3920));
  nor2 g03727(.a(new_n2660), .b(new_n257), .O(new_n3921));
  inv1 g03728(.a(new_n3921), .O(new_n3922));
  nor2 g03729(.a(new_n2433), .b(new_n322), .O(new_n3923));
  nor2 g03730(.a(new_n2506), .b(new_n295), .O(new_n3924));
  nor2 g03731(.a(new_n3924), .b(new_n3923), .O(new_n3925));
  nor2 g03732(.a(new_n3683), .b(new_n3674), .O(new_n3926));
  nor2 g03733(.a(new_n3926), .b(new_n3925), .O(new_n3927));
  nor2 g03734(.a(new_n3927), .b(new_n3922), .O(new_n3928));
  inv1 g03735(.a(new_n3927), .O(new_n3929));
  nor2 g03736(.a(new_n3929), .b(new_n3921), .O(new_n3930));
  nor2 g03737(.a(new_n3930), .b(new_n3928), .O(new_n3931));
  inv1 g03738(.a(new_n3931), .O(new_n3932));
  nor2 g03739(.a(new_n3533), .b(new_n196), .O(new_n3933));
  nor2 g03740(.a(new_n1647), .b(new_n613), .O(new_n3934));
  nor2 g03741(.a(new_n3934), .b(new_n3741), .O(new_n3935));
  nor2 g03742(.a(new_n1736), .b(new_n613), .O(new_n3936));
  inv1 g03743(.a(new_n3936), .O(new_n3937));
  nor2 g03744(.a(new_n3937), .b(new_n3440), .O(new_n3938));
  nor2 g03745(.a(new_n3938), .b(new_n3935), .O(new_n3939));
  inv1 g03746(.a(new_n3939), .O(new_n3940));
  nor2 g03747(.a(new_n3940), .b(new_n3933), .O(new_n3941));
  inv1 g03748(.a(new_n3933), .O(new_n3942));
  nor2 g03749(.a(new_n3939), .b(new_n3942), .O(new_n3943));
  nor2 g03750(.a(new_n3943), .b(new_n3941), .O(new_n3944));
  nor2 g03751(.a(new_n2826), .b(new_n229), .O(new_n3945));
  nor2 g03752(.a(new_n2184), .b(new_n363), .O(new_n3946));
  nor2 g03753(.a(new_n3946), .b(new_n3945), .O(new_n3947));
  inv1 g03754(.a(new_n3011), .O(new_n3948));
  nor2 g03755(.a(new_n3948), .b(new_n2831), .O(new_n3949));
  nor2 g03756(.a(new_n3949), .b(new_n3947), .O(new_n3950));
  nor2 g03757(.a(new_n3950), .b(new_n3661), .O(new_n3951));
  inv1 g03758(.a(new_n3950), .O(new_n3952));
  nor2 g03759(.a(new_n3952), .b(new_n3660), .O(new_n3953));
  nor2 g03760(.a(new_n3953), .b(new_n3951), .O(new_n3954));
  nor2 g03761(.a(new_n3954), .b(new_n3944), .O(new_n3955));
  inv1 g03762(.a(new_n3944), .O(new_n3956));
  inv1 g03763(.a(new_n3954), .O(new_n3957));
  nor2 g03764(.a(new_n3957), .b(new_n3956), .O(new_n3958));
  nor2 g03765(.a(new_n3958), .b(new_n3955), .O(new_n3959));
  nor2 g03766(.a(new_n3959), .b(new_n3932), .O(new_n3960));
  inv1 g03767(.a(new_n3959), .O(new_n3961));
  nor2 g03768(.a(new_n3961), .b(new_n3931), .O(new_n3962));
  nor2 g03769(.a(new_n3962), .b(new_n3960), .O(new_n3963));
  inv1 g03770(.a(new_n3963), .O(new_n3964));
  nor2 g03771(.a(new_n3964), .b(new_n3920), .O(new_n3965));
  nor2 g03772(.a(new_n3963), .b(new_n3919), .O(new_n3966));
  nor2 g03773(.a(new_n3966), .b(new_n3965), .O(new_n3967));
  inv1 g03774(.a(new_n3967), .O(new_n3968));
  nor2 g03775(.a(new_n3968), .b(new_n3859), .O(new_n3969));
  nor2 g03776(.a(new_n3967), .b(new_n3858), .O(new_n3970));
  nor2 g03777(.a(new_n3970), .b(new_n3969), .O(new_n3971));
  inv1 g03778(.a(new_n3971), .O(new_n3972));
  nor2 g03779(.a(new_n3972), .b(new_n3815), .O(new_n3973));
  nor2 g03780(.a(new_n3971), .b(new_n3814), .O(new_n3974));
  nor2 g03781(.a(new_n3974), .b(new_n3973), .O(new_n3975));
  nor2 g03782(.a(new_n3975), .b(new_n3783), .O(new_n3976));
  inv1 g03783(.a(new_n3975), .O(new_n3977));
  nor2 g03784(.a(new_n3977), .b(new_n3782), .O(new_n3978));
  nor2 g03785(.a(new_n3978), .b(new_n3976), .O(new_n3979));
  nor2 g03786(.a(new_n3777), .b(new_n3771), .O(new_n3980));
  inv1 g03787(.a(new_n3980), .O(new_n3981));
  nor2 g03788(.a(new_n3981), .b(new_n3979), .O(new_n3982));
  inv1 g03789(.a(new_n3979), .O(new_n3983));
  nor2 g03790(.a(new_n3980), .b(new_n3983), .O(new_n3984));
  nor2 g03791(.a(new_n3984), .b(new_n3982), .O(new_n3985));
  inv1 g03792(.a(new_n3985), .O(\asquared[37] ));
  nor2 g03793(.a(new_n3973), .b(new_n3811), .O(new_n3987));
  nor2 g03794(.a(new_n3806), .b(new_n3802), .O(new_n3988));
  nor2 g03795(.a(new_n3904), .b(new_n3897), .O(new_n3989));
  nor2 g03796(.a(new_n3891), .b(new_n3884), .O(new_n3990));
  nor2 g03797(.a(new_n3990), .b(new_n3989), .O(new_n3991));
  inv1 g03798(.a(new_n3989), .O(new_n3992));
  inv1 g03799(.a(new_n3990), .O(new_n3993));
  nor2 g03800(.a(new_n3993), .b(new_n3992), .O(new_n3994));
  nor2 g03801(.a(new_n3994), .b(new_n3991), .O(new_n3995));
  nor2 g03802(.a(new_n3941), .b(new_n3935), .O(new_n3996));
  nor2 g03803(.a(new_n3996), .b(new_n3995), .O(new_n3997));
  inv1 g03804(.a(new_n3995), .O(new_n3998));
  inv1 g03805(.a(new_n3996), .O(new_n3999));
  nor2 g03806(.a(new_n3999), .b(new_n3998), .O(new_n4000));
  nor2 g03807(.a(new_n4000), .b(new_n3997), .O(new_n4001));
  inv1 g03808(.a(new_n4001), .O(new_n4002));
  nor2 g03809(.a(new_n3912), .b(new_n3906), .O(new_n4003));
  nor2 g03810(.a(new_n4003), .b(new_n4002), .O(new_n4004));
  inv1 g03811(.a(new_n4003), .O(new_n4005));
  nor2 g03812(.a(new_n4005), .b(new_n4001), .O(new_n4006));
  nor2 g03813(.a(new_n4006), .b(new_n4004), .O(new_n4007));
  inv1 g03814(.a(new_n4007), .O(new_n4008));
  nor2 g03815(.a(new_n3877), .b(new_n3873), .O(new_n4009));
  inv1 g03816(.a(new_n4009), .O(new_n4010));
  nor2 g03817(.a(new_n3953), .b(new_n3947), .O(new_n4011));
  nor2 g03818(.a(new_n4011), .b(new_n4010), .O(new_n4012));
  inv1 g03819(.a(new_n4011), .O(new_n4013));
  nor2 g03820(.a(new_n4013), .b(new_n4009), .O(new_n4014));
  nor2 g03821(.a(new_n4014), .b(new_n4012), .O(new_n4015));
  inv1 g03822(.a(new_n4015), .O(new_n4016));
  nor2 g03823(.a(new_n1647), .b(new_n699), .O(new_n4017));
  nor2 g03824(.a(new_n1493), .b(new_n800), .O(new_n4018));
  nor2 g03825(.a(new_n4018), .b(new_n4017), .O(new_n4019));
  nor2 g03826(.a(new_n1647), .b(new_n800), .O(new_n4020));
  inv1 g03827(.a(new_n4020), .O(new_n4021));
  nor2 g03828(.a(new_n4021), .b(new_n3882), .O(new_n4022));
  nor2 g03829(.a(new_n4022), .b(new_n4019), .O(new_n4023));
  nor2 g03830(.a(new_n4023), .b(new_n3937), .O(new_n4024));
  inv1 g03831(.a(new_n4023), .O(new_n4025));
  nor2 g03832(.a(new_n4025), .b(new_n3936), .O(new_n4026));
  nor2 g03833(.a(new_n4026), .b(new_n4024), .O(new_n4027));
  nor2 g03834(.a(new_n4027), .b(new_n4016), .O(new_n4028));
  inv1 g03835(.a(new_n4027), .O(new_n4029));
  nor2 g03836(.a(new_n4029), .b(new_n4015), .O(new_n4030));
  nor2 g03837(.a(new_n4030), .b(new_n4028), .O(new_n4031));
  inv1 g03838(.a(new_n4031), .O(new_n4032));
  nor2 g03839(.a(new_n4032), .b(new_n4008), .O(new_n4033));
  nor2 g03840(.a(new_n4031), .b(new_n4007), .O(new_n4034));
  nor2 g03841(.a(new_n4034), .b(new_n4033), .O(new_n4035));
  inv1 g03842(.a(new_n4035), .O(new_n4036));
  nor2 g03843(.a(new_n4036), .b(new_n3988), .O(new_n4037));
  inv1 g03844(.a(new_n3988), .O(new_n4038));
  nor2 g03845(.a(new_n4035), .b(new_n4038), .O(new_n4039));
  nor2 g03846(.a(new_n4039), .b(new_n4037), .O(new_n4040));
  inv1 g03847(.a(new_n4040), .O(new_n4041));
  nor2 g03848(.a(new_n3842), .b(new_n3836), .O(new_n4042));
  inv1 g03849(.a(new_n4042), .O(new_n4043));
  nor2 g03850(.a(new_n2121), .b(new_n502), .O(new_n4044));
  nor2 g03851(.a(new_n3057), .b(new_n229), .O(new_n4045));
  nor2 g03852(.a(new_n2184), .b(new_n438), .O(new_n4046));
  nor2 g03853(.a(new_n4046), .b(new_n4045), .O(new_n4047));
  nor2 g03854(.a(new_n3057), .b(new_n438), .O(new_n4048));
  inv1 g03855(.a(new_n4048), .O(new_n4049));
  nor2 g03856(.a(new_n4049), .b(new_n3948), .O(new_n4050));
  nor2 g03857(.a(new_n4050), .b(new_n4047), .O(new_n4051));
  inv1 g03858(.a(new_n4051), .O(new_n4052));
  nor2 g03859(.a(new_n4052), .b(new_n4044), .O(new_n4053));
  inv1 g03860(.a(new_n4044), .O(new_n4054));
  nor2 g03861(.a(new_n4051), .b(new_n4054), .O(new_n4055));
  nor2 g03862(.a(new_n4055), .b(new_n4053), .O(new_n4056));
  nor2 g03863(.a(new_n1199), .b(new_n1086), .O(new_n4057));
  nor2 g03864(.a(new_n1297), .b(new_n941), .O(new_n4058));
  nor2 g03865(.a(new_n4058), .b(new_n4057), .O(new_n4059));
  nor2 g03866(.a(new_n1297), .b(new_n1086), .O(new_n4060));
  inv1 g03867(.a(new_n4060), .O(new_n4061));
  nor2 g03868(.a(new_n4061), .b(new_n3864), .O(new_n4062));
  nor2 g03869(.a(new_n4062), .b(new_n4059), .O(new_n4063));
  nor2 g03870(.a(new_n4063), .b(new_n3674), .O(new_n4064));
  inv1 g03871(.a(new_n4063), .O(new_n4065));
  nor2 g03872(.a(new_n4065), .b(new_n3673), .O(new_n4066));
  nor2 g03873(.a(new_n4066), .b(new_n4064), .O(new_n4067));
  nor2 g03874(.a(new_n4067), .b(new_n4056), .O(new_n4068));
  inv1 g03875(.a(new_n4056), .O(new_n4069));
  inv1 g03876(.a(new_n4067), .O(new_n4070));
  nor2 g03877(.a(new_n4070), .b(new_n4069), .O(new_n4071));
  nor2 g03878(.a(new_n4071), .b(new_n4068), .O(new_n4072));
  nor2 g03879(.a(new_n4072), .b(new_n4043), .O(new_n4073));
  inv1 g03880(.a(new_n4072), .O(new_n4074));
  nor2 g03881(.a(new_n4074), .b(new_n4042), .O(new_n4075));
  nor2 g03882(.a(new_n4075), .b(new_n4073), .O(new_n4076));
  nor2 g03883(.a(new_n3796), .b(new_n3790), .O(new_n4077));
  inv1 g03884(.a(new_n4077), .O(new_n4078));
  nor2 g03885(.a(new_n4078), .b(new_n4076), .O(new_n4079));
  inv1 g03886(.a(new_n4076), .O(new_n4080));
  nor2 g03887(.a(new_n4077), .b(new_n4080), .O(new_n4081));
  nor2 g03888(.a(new_n4081), .b(new_n4079), .O(new_n4082));
  nor2 g03889(.a(new_n3533), .b(new_n203), .O(new_n4083));
  nor2 g03890(.a(new_n4083), .b(new_n3727), .O(new_n4084));
  nor2 g03891(.a(new_n3722), .b(new_n203), .O(new_n4085));
  inv1 g03892(.a(new_n4085), .O(new_n4086));
  nor2 g03893(.a(new_n4086), .b(new_n3942), .O(new_n4087));
  nor2 g03894(.a(new_n4087), .b(new_n4084), .O(new_n4088));
  nor2 g03895(.a(new_n4088), .b(new_n3886), .O(new_n4089));
  inv1 g03896(.a(new_n4088), .O(new_n4090));
  nor2 g03897(.a(new_n4090), .b(new_n3885), .O(new_n4091));
  nor2 g03898(.a(new_n4091), .b(new_n4089), .O(new_n4092));
  inv1 g03899(.a(\a[37] ), .O(new_n4093));
  nor2 g03900(.a(new_n4093), .b(new_n198), .O(new_n4094));
  inv1 g03901(.a(new_n4094), .O(new_n4095));
  nor2 g03902(.a(new_n1903), .b(new_n569), .O(new_n4096));
  nor2 g03903(.a(new_n3231), .b(new_n214), .O(new_n4097));
  nor2 g03904(.a(new_n4097), .b(new_n4096), .O(new_n4098));
  nor2 g03905(.a(new_n3231), .b(new_n569), .O(new_n4099));
  inv1 g03906(.a(new_n4099), .O(new_n4100));
  nor2 g03907(.a(new_n4100), .b(new_n2339), .O(new_n4101));
  nor2 g03908(.a(new_n4101), .b(new_n4098), .O(new_n4102));
  nor2 g03909(.a(new_n4102), .b(new_n4095), .O(new_n4103));
  inv1 g03910(.a(new_n4102), .O(new_n4104));
  nor2 g03911(.a(new_n4104), .b(new_n4094), .O(new_n4105));
  nor2 g03912(.a(new_n4105), .b(new_n4103), .O(new_n4106));
  nor2 g03913(.a(new_n4106), .b(new_n4092), .O(new_n4107));
  inv1 g03914(.a(new_n4092), .O(new_n4108));
  inv1 g03915(.a(new_n4106), .O(new_n4109));
  nor2 g03916(.a(new_n4109), .b(new_n4108), .O(new_n4110));
  nor2 g03917(.a(new_n4110), .b(new_n4107), .O(new_n4111));
  inv1 g03918(.a(new_n4111), .O(new_n4112));
  nor2 g03919(.a(new_n2433), .b(new_n363), .O(new_n4113));
  inv1 g03920(.a(new_n4113), .O(new_n4114));
  nor2 g03921(.a(new_n2826), .b(new_n257), .O(new_n4115));
  nor2 g03922(.a(new_n2660), .b(new_n295), .O(new_n4116));
  nor2 g03923(.a(new_n4116), .b(new_n4115), .O(new_n4117));
  nor2 g03924(.a(new_n2826), .b(new_n295), .O(new_n4118));
  inv1 g03925(.a(new_n4118), .O(new_n4119));
  nor2 g03926(.a(new_n4119), .b(new_n3922), .O(new_n4120));
  nor2 g03927(.a(new_n4120), .b(new_n4117), .O(new_n4121));
  nor2 g03928(.a(new_n4121), .b(new_n4114), .O(new_n4122));
  inv1 g03929(.a(new_n4121), .O(new_n4123));
  nor2 g03930(.a(new_n4123), .b(new_n4113), .O(new_n4124));
  nor2 g03931(.a(new_n4124), .b(new_n4122), .O(new_n4125));
  nor2 g03932(.a(new_n4125), .b(new_n4112), .O(new_n4126));
  inv1 g03933(.a(new_n4125), .O(new_n4127));
  nor2 g03934(.a(new_n4127), .b(new_n4111), .O(new_n4128));
  nor2 g03935(.a(new_n4128), .b(new_n4126), .O(new_n4129));
  nor2 g03936(.a(new_n4129), .b(new_n4082), .O(new_n4130));
  inv1 g03937(.a(new_n4082), .O(new_n4131));
  inv1 g03938(.a(new_n4129), .O(new_n4132));
  nor2 g03939(.a(new_n4132), .b(new_n4131), .O(new_n4133));
  nor2 g03940(.a(new_n4133), .b(new_n4130), .O(new_n4134));
  inv1 g03941(.a(new_n4134), .O(new_n4135));
  nor2 g03942(.a(new_n4135), .b(new_n4041), .O(new_n4136));
  nor2 g03943(.a(new_n4134), .b(new_n4040), .O(new_n4137));
  nor2 g03944(.a(new_n4137), .b(new_n4136), .O(new_n4138));
  inv1 g03945(.a(new_n4138), .O(new_n4139));
  nor2 g03946(.a(new_n3969), .b(new_n3855), .O(new_n4140));
  nor2 g03947(.a(new_n3851), .b(new_n3848), .O(new_n4141));
  nor2 g03948(.a(new_n3828), .b(new_n3822), .O(new_n4142));
  inv1 g03949(.a(new_n3866), .O(new_n4143));
  nor2 g03950(.a(new_n4143), .b(\a[36] ), .O(new_n4144));
  nor2 g03951(.a(new_n1276), .b(new_n3870), .O(new_n4145));
  nor2 g03952(.a(new_n3870), .b(new_n194), .O(new_n4146));
  nor2 g03953(.a(new_n4146), .b(\a[19] ), .O(new_n4147));
  nor2 g03954(.a(new_n4147), .b(new_n4145), .O(new_n4148));
  nor2 g03955(.a(new_n4148), .b(new_n3866), .O(new_n4149));
  nor2 g03956(.a(new_n4149), .b(new_n4144), .O(new_n4150));
  inv1 g03957(.a(new_n4150), .O(new_n4151));
  nor2 g03958(.a(new_n3930), .b(new_n3925), .O(new_n4152));
  inv1 g03959(.a(new_n4152), .O(new_n4153));
  nor2 g03960(.a(new_n4153), .b(new_n4151), .O(new_n4154));
  nor2 g03961(.a(new_n4152), .b(new_n4150), .O(new_n4155));
  nor2 g03962(.a(new_n4155), .b(new_n4154), .O(new_n4156));
  inv1 g03963(.a(new_n4156), .O(new_n4157));
  nor2 g03964(.a(new_n4157), .b(new_n4142), .O(new_n4158));
  inv1 g03965(.a(new_n4142), .O(new_n4159));
  nor2 g03966(.a(new_n4156), .b(new_n4159), .O(new_n4160));
  nor2 g03967(.a(new_n4160), .b(new_n4158), .O(new_n4161));
  inv1 g03968(.a(new_n4161), .O(new_n4162));
  nor2 g03969(.a(new_n3962), .b(new_n3955), .O(new_n4163));
  nor2 g03970(.a(new_n4163), .b(new_n4162), .O(new_n4164));
  inv1 g03971(.a(new_n4163), .O(new_n4165));
  nor2 g03972(.a(new_n4165), .b(new_n4161), .O(new_n4166));
  nor2 g03973(.a(new_n4166), .b(new_n4164), .O(new_n4167));
  inv1 g03974(.a(new_n4167), .O(new_n4168));
  nor2 g03975(.a(new_n4168), .b(new_n4141), .O(new_n4169));
  inv1 g03976(.a(new_n4141), .O(new_n4170));
  nor2 g03977(.a(new_n4167), .b(new_n4170), .O(new_n4171));
  nor2 g03978(.a(new_n4171), .b(new_n4169), .O(new_n4172));
  inv1 g03979(.a(new_n4172), .O(new_n4173));
  nor2 g03980(.a(new_n3965), .b(new_n3916), .O(new_n4174));
  nor2 g03981(.a(new_n4174), .b(new_n4173), .O(new_n4175));
  inv1 g03982(.a(new_n4174), .O(new_n4176));
  nor2 g03983(.a(new_n4176), .b(new_n4172), .O(new_n4177));
  nor2 g03984(.a(new_n4177), .b(new_n4175), .O(new_n4178));
  inv1 g03985(.a(new_n4178), .O(new_n4179));
  nor2 g03986(.a(new_n4179), .b(new_n4140), .O(new_n4180));
  inv1 g03987(.a(new_n4140), .O(new_n4181));
  nor2 g03988(.a(new_n4178), .b(new_n4181), .O(new_n4182));
  nor2 g03989(.a(new_n4182), .b(new_n4180), .O(new_n4183));
  inv1 g03990(.a(new_n4183), .O(new_n4184));
  nor2 g03991(.a(new_n4184), .b(new_n4139), .O(new_n4185));
  nor2 g03992(.a(new_n4183), .b(new_n4138), .O(new_n4186));
  nor2 g03993(.a(new_n4186), .b(new_n4185), .O(new_n4187));
  inv1 g03994(.a(new_n4187), .O(new_n4188));
  nor2 g03995(.a(new_n4188), .b(new_n3987), .O(new_n4189));
  inv1 g03996(.a(new_n3987), .O(new_n4190));
  nor2 g03997(.a(new_n4187), .b(new_n4190), .O(new_n4191));
  nor2 g03998(.a(new_n4191), .b(new_n4189), .O(new_n4192));
  inv1 g03999(.a(new_n4192), .O(new_n4193));
  nor2 g04000(.a(new_n3984), .b(new_n3976), .O(new_n4194));
  nor2 g04001(.a(new_n4194), .b(new_n4193), .O(new_n4195));
  inv1 g04002(.a(new_n4194), .O(new_n4196));
  nor2 g04003(.a(new_n4196), .b(new_n4192), .O(new_n4197));
  nor2 g04004(.a(new_n4197), .b(new_n4195), .O(new_n4198));
  inv1 g04005(.a(new_n4198), .O(\asquared[38] ));
  nor2 g04006(.a(new_n4185), .b(new_n4180), .O(new_n4200));
  nor2 g04007(.a(new_n4136), .b(new_n4037), .O(new_n4201));
  inv1 g04008(.a(new_n4201), .O(new_n4202));
  nor2 g04009(.a(new_n4105), .b(new_n4098), .O(new_n4203));
  nor2 g04010(.a(new_n4091), .b(new_n4084), .O(new_n4204));
  nor2 g04011(.a(new_n4204), .b(new_n4203), .O(new_n4205));
  inv1 g04012(.a(new_n4203), .O(new_n4206));
  inv1 g04013(.a(new_n4204), .O(new_n4207));
  nor2 g04014(.a(new_n4207), .b(new_n4206), .O(new_n4208));
  nor2 g04015(.a(new_n4208), .b(new_n4205), .O(new_n4209));
  nor2 g04016(.a(new_n4026), .b(new_n4019), .O(new_n4210));
  nor2 g04017(.a(new_n4210), .b(new_n4209), .O(new_n4211));
  inv1 g04018(.a(new_n4209), .O(new_n4212));
  inv1 g04019(.a(new_n4210), .O(new_n4213));
  nor2 g04020(.a(new_n4213), .b(new_n4212), .O(new_n4214));
  nor2 g04021(.a(new_n4214), .b(new_n4211), .O(new_n4215));
  nor2 g04022(.a(new_n4075), .b(new_n4068), .O(new_n4216));
  inv1 g04023(.a(new_n4216), .O(new_n4217));
  nor2 g04024(.a(new_n4217), .b(new_n4215), .O(new_n4218));
  inv1 g04025(.a(new_n4215), .O(new_n4219));
  nor2 g04026(.a(new_n4216), .b(new_n4219), .O(new_n4220));
  nor2 g04027(.a(new_n4220), .b(new_n4218), .O(new_n4221));
  inv1 g04028(.a(new_n4221), .O(new_n4222));
  nor2 g04029(.a(new_n2506), .b(new_n363), .O(new_n4223));
  inv1 g04030(.a(new_n4223), .O(new_n4224));
  nor2 g04031(.a(new_n2660), .b(new_n322), .O(new_n4225));
  nor2 g04032(.a(new_n4225), .b(new_n4118), .O(new_n4226));
  inv1 g04033(.a(new_n4116), .O(new_n4227));
  nor2 g04034(.a(new_n2826), .b(new_n322), .O(new_n4228));
  inv1 g04035(.a(new_n4228), .O(new_n4229));
  nor2 g04036(.a(new_n4229), .b(new_n4227), .O(new_n4230));
  nor2 g04037(.a(new_n4230), .b(new_n4226), .O(new_n4231));
  nor2 g04038(.a(new_n4231), .b(new_n4224), .O(new_n4232));
  inv1 g04039(.a(new_n4231), .O(new_n4233));
  nor2 g04040(.a(new_n4233), .b(new_n4223), .O(new_n4234));
  nor2 g04041(.a(new_n4234), .b(new_n4232), .O(new_n4235));
  nor2 g04042(.a(new_n1493), .b(new_n847), .O(new_n4236));
  nor2 g04043(.a(new_n1425), .b(new_n941), .O(new_n4237));
  nor2 g04044(.a(new_n4237), .b(new_n4236), .O(new_n4238));
  nor2 g04045(.a(new_n1493), .b(new_n941), .O(new_n4239));
  inv1 g04046(.a(new_n4239), .O(new_n4240));
  nor2 g04047(.a(new_n4240), .b(new_n3886), .O(new_n4241));
  nor2 g04048(.a(new_n4241), .b(new_n4238), .O(new_n4242));
  nor2 g04049(.a(new_n4242), .b(new_n4021), .O(new_n4243));
  inv1 g04050(.a(new_n4242), .O(new_n4244));
  nor2 g04051(.a(new_n4244), .b(new_n4020), .O(new_n4245));
  nor2 g04052(.a(new_n4245), .b(new_n4243), .O(new_n4246));
  nor2 g04053(.a(new_n3231), .b(new_n229), .O(new_n4247));
  inv1 g04054(.a(new_n4247), .O(new_n4248));
  nor2 g04055(.a(new_n2433), .b(new_n438), .O(new_n4249));
  nor2 g04056(.a(new_n3057), .b(new_n257), .O(new_n4250));
  nor2 g04057(.a(new_n4250), .b(new_n4249), .O(new_n4251));
  inv1 g04058(.a(new_n4249), .O(new_n4252));
  inv1 g04059(.a(new_n4250), .O(new_n4253));
  nor2 g04060(.a(new_n4253), .b(new_n4252), .O(new_n4254));
  nor2 g04061(.a(new_n4254), .b(new_n4251), .O(new_n4255));
  nor2 g04062(.a(new_n4255), .b(new_n4248), .O(new_n4256));
  inv1 g04063(.a(new_n4255), .O(new_n4257));
  nor2 g04064(.a(new_n4257), .b(new_n4247), .O(new_n4258));
  nor2 g04065(.a(new_n4258), .b(new_n4256), .O(new_n4259));
  nor2 g04066(.a(new_n4259), .b(new_n4246), .O(new_n4260));
  inv1 g04067(.a(new_n4246), .O(new_n4261));
  inv1 g04068(.a(new_n4259), .O(new_n4262));
  nor2 g04069(.a(new_n4262), .b(new_n4261), .O(new_n4263));
  nor2 g04070(.a(new_n4263), .b(new_n4260), .O(new_n4264));
  inv1 g04071(.a(new_n4264), .O(new_n4265));
  nor2 g04072(.a(new_n4265), .b(new_n4235), .O(new_n4266));
  inv1 g04073(.a(new_n4235), .O(new_n4267));
  nor2 g04074(.a(new_n4264), .b(new_n4267), .O(new_n4268));
  nor2 g04075(.a(new_n4268), .b(new_n4266), .O(new_n4269));
  inv1 g04076(.a(new_n4269), .O(new_n4270));
  nor2 g04077(.a(new_n4270), .b(new_n4222), .O(new_n4271));
  nor2 g04078(.a(new_n4269), .b(new_n4221), .O(new_n4272));
  nor2 g04079(.a(new_n4272), .b(new_n4271), .O(new_n4273));
  inv1 g04080(.a(new_n4273), .O(new_n4274));
  nor2 g04081(.a(new_n4133), .b(new_n4081), .O(new_n4275));
  nor2 g04082(.a(new_n4033), .b(new_n4004), .O(new_n4276));
  nor2 g04083(.a(new_n4276), .b(new_n4275), .O(new_n4277));
  inv1 g04084(.a(new_n4275), .O(new_n4278));
  inv1 g04085(.a(new_n4276), .O(new_n4279));
  nor2 g04086(.a(new_n4279), .b(new_n4278), .O(new_n4280));
  nor2 g04087(.a(new_n4280), .b(new_n4277), .O(new_n4281));
  inv1 g04088(.a(new_n4281), .O(new_n4282));
  nor2 g04089(.a(new_n4282), .b(new_n4274), .O(new_n4283));
  nor2 g04090(.a(new_n4281), .b(new_n4273), .O(new_n4284));
  nor2 g04091(.a(new_n4284), .b(new_n4283), .O(new_n4285));
  nor2 g04092(.a(new_n4285), .b(new_n4202), .O(new_n4286));
  inv1 g04093(.a(new_n4285), .O(new_n4287));
  nor2 g04094(.a(new_n4287), .b(new_n4201), .O(new_n4288));
  nor2 g04095(.a(new_n4288), .b(new_n4286), .O(new_n4289));
  nor2 g04096(.a(new_n4175), .b(new_n4169), .O(new_n4290));
  inv1 g04097(.a(new_n4290), .O(new_n4291));
  nor2 g04098(.a(new_n4126), .b(new_n4107), .O(new_n4292));
  inv1 g04099(.a(new_n4292), .O(new_n4293));
  nor2 g04100(.a(new_n4028), .b(new_n4014), .O(new_n4294));
  inv1 g04101(.a(new_n4294), .O(new_n4295));
  nor2 g04102(.a(new_n4295), .b(new_n4293), .O(new_n4296));
  nor2 g04103(.a(new_n4294), .b(new_n4292), .O(new_n4297));
  nor2 g04104(.a(new_n4297), .b(new_n4296), .O(new_n4298));
  inv1 g04105(.a(new_n4298), .O(new_n4299));
  nor2 g04106(.a(new_n4093), .b(new_n194), .O(new_n4300));
  nor2 g04107(.a(new_n4300), .b(new_n4060), .O(new_n4301));
  inv1 g04108(.a(new_n4300), .O(new_n4302));
  nor2 g04109(.a(new_n4302), .b(new_n4061), .O(new_n4303));
  nor2 g04110(.a(new_n4303), .b(new_n4301), .O(new_n4304));
  nor2 g04111(.a(new_n4066), .b(new_n4059), .O(new_n4305));
  nor2 g04112(.a(new_n4305), .b(new_n4304), .O(new_n4306));
  inv1 g04113(.a(new_n4304), .O(new_n4307));
  inv1 g04114(.a(new_n4305), .O(new_n4308));
  nor2 g04115(.a(new_n4308), .b(new_n4307), .O(new_n4309));
  nor2 g04116(.a(new_n4309), .b(new_n4306), .O(new_n4310));
  inv1 g04117(.a(new_n4310), .O(new_n4311));
  nor2 g04118(.a(new_n4124), .b(new_n4117), .O(new_n4312));
  inv1 g04119(.a(new_n4312), .O(new_n4313));
  nor2 g04120(.a(new_n4313), .b(new_n4311), .O(new_n4314));
  nor2 g04121(.a(new_n4312), .b(new_n4310), .O(new_n4315));
  nor2 g04122(.a(new_n4315), .b(new_n4314), .O(new_n4316));
  inv1 g04123(.a(new_n4316), .O(new_n4317));
  nor2 g04124(.a(new_n4317), .b(new_n4299), .O(new_n4318));
  nor2 g04125(.a(new_n4316), .b(new_n4298), .O(new_n4319));
  nor2 g04126(.a(new_n4319), .b(new_n4318), .O(new_n4320));
  nor2 g04127(.a(new_n4320), .b(new_n4291), .O(new_n4321));
  inv1 g04128(.a(new_n4320), .O(new_n4322));
  nor2 g04129(.a(new_n4322), .b(new_n4290), .O(new_n4323));
  nor2 g04130(.a(new_n4323), .b(new_n4321), .O(new_n4324));
  inv1 g04131(.a(new_n4324), .O(new_n4325));
  nor2 g04132(.a(new_n4000), .b(new_n3994), .O(new_n4326));
  inv1 g04133(.a(new_n4326), .O(new_n4327));
  nor2 g04134(.a(new_n4154), .b(new_n4144), .O(new_n4328));
  nor2 g04135(.a(new_n2121), .b(new_n569), .O(new_n4329));
  inv1 g04136(.a(new_n4329), .O(new_n4330));
  nor2 g04137(.a(new_n3533), .b(new_n214), .O(new_n4331));
  nor2 g04138(.a(new_n2184), .b(new_n502), .O(new_n4332));
  nor2 g04139(.a(new_n4332), .b(new_n4331), .O(new_n4333));
  nor2 g04140(.a(new_n3533), .b(new_n502), .O(new_n4334));
  inv1 g04141(.a(new_n4334), .O(new_n4335));
  nor2 g04142(.a(new_n4335), .b(new_n3013), .O(new_n4336));
  nor2 g04143(.a(new_n4336), .b(new_n4333), .O(new_n4337));
  nor2 g04144(.a(new_n4337), .b(new_n4330), .O(new_n4338));
  inv1 g04145(.a(new_n4337), .O(new_n4339));
  nor2 g04146(.a(new_n4339), .b(new_n4329), .O(new_n4340));
  nor2 g04147(.a(new_n4340), .b(new_n4338), .O(new_n4341));
  nor2 g04148(.a(new_n4341), .b(new_n4328), .O(new_n4342));
  inv1 g04149(.a(new_n4328), .O(new_n4343));
  inv1 g04150(.a(new_n4341), .O(new_n4344));
  nor2 g04151(.a(new_n4344), .b(new_n4343), .O(new_n4345));
  nor2 g04152(.a(new_n4345), .b(new_n4342), .O(new_n4346));
  nor2 g04153(.a(new_n4346), .b(new_n4327), .O(new_n4347));
  inv1 g04154(.a(new_n4346), .O(new_n4348));
  nor2 g04155(.a(new_n4348), .b(new_n4326), .O(new_n4349));
  nor2 g04156(.a(new_n4349), .b(new_n4347), .O(new_n4350));
  inv1 g04157(.a(new_n4350), .O(new_n4351));
  nor2 g04158(.a(new_n4164), .b(new_n4158), .O(new_n4352));
  inv1 g04159(.a(new_n4352), .O(new_n4353));
  nor2 g04160(.a(new_n1903), .b(new_n613), .O(new_n4354));
  nor2 g04161(.a(new_n1736), .b(new_n699), .O(new_n4355));
  nor2 g04162(.a(new_n4355), .b(new_n4354), .O(new_n4356));
  nor2 g04163(.a(new_n1903), .b(new_n699), .O(new_n4357));
  inv1 g04164(.a(new_n4357), .O(new_n4358));
  nor2 g04165(.a(new_n4358), .b(new_n3937), .O(new_n4359));
  nor2 g04166(.a(new_n4359), .b(new_n4356), .O(new_n4360));
  nor2 g04167(.a(new_n4360), .b(new_n4086), .O(new_n4361));
  inv1 g04168(.a(new_n4360), .O(new_n4362));
  nor2 g04169(.a(new_n4362), .b(new_n4085), .O(new_n4363));
  nor2 g04170(.a(new_n4363), .b(new_n4361), .O(new_n4364));
  inv1 g04171(.a(new_n4145), .O(new_n4365));
  inv1 g04172(.a(\a[38] ), .O(new_n4366));
  nor2 g04173(.a(new_n4366), .b(new_n198), .O(new_n4367));
  nor2 g04174(.a(new_n3870), .b(new_n196), .O(new_n4368));
  nor2 g04175(.a(new_n4368), .b(new_n4367), .O(new_n4369));
  nor2 g04176(.a(new_n4366), .b(new_n196), .O(new_n4370));
  inv1 g04177(.a(new_n4370), .O(new_n4371));
  nor2 g04178(.a(new_n4371), .b(new_n3872), .O(new_n4372));
  nor2 g04179(.a(new_n4372), .b(new_n4369), .O(new_n4373));
  nor2 g04180(.a(new_n4373), .b(new_n4365), .O(new_n4374));
  inv1 g04181(.a(new_n4373), .O(new_n4375));
  nor2 g04182(.a(new_n4375), .b(new_n4145), .O(new_n4376));
  nor2 g04183(.a(new_n4376), .b(new_n4374), .O(new_n4377));
  nor2 g04184(.a(new_n4053), .b(new_n4047), .O(new_n4378));
  inv1 g04185(.a(new_n4378), .O(new_n4379));
  nor2 g04186(.a(new_n4379), .b(new_n4377), .O(new_n4380));
  inv1 g04187(.a(new_n4377), .O(new_n4381));
  nor2 g04188(.a(new_n4378), .b(new_n4381), .O(new_n4382));
  nor2 g04189(.a(new_n4382), .b(new_n4380), .O(new_n4383));
  inv1 g04190(.a(new_n4383), .O(new_n4384));
  nor2 g04191(.a(new_n4384), .b(new_n4364), .O(new_n4385));
  inv1 g04192(.a(new_n4364), .O(new_n4386));
  nor2 g04193(.a(new_n4383), .b(new_n4386), .O(new_n4387));
  nor2 g04194(.a(new_n4387), .b(new_n4385), .O(new_n4388));
  nor2 g04195(.a(new_n4388), .b(new_n4353), .O(new_n4389));
  inv1 g04196(.a(new_n4388), .O(new_n4390));
  nor2 g04197(.a(new_n4390), .b(new_n4352), .O(new_n4391));
  nor2 g04198(.a(new_n4391), .b(new_n4389), .O(new_n4392));
  inv1 g04199(.a(new_n4392), .O(new_n4393));
  nor2 g04200(.a(new_n4393), .b(new_n4351), .O(new_n4394));
  nor2 g04201(.a(new_n4392), .b(new_n4350), .O(new_n4395));
  nor2 g04202(.a(new_n4395), .b(new_n4394), .O(new_n4396));
  inv1 g04203(.a(new_n4396), .O(new_n4397));
  nor2 g04204(.a(new_n4397), .b(new_n4325), .O(new_n4398));
  nor2 g04205(.a(new_n4396), .b(new_n4324), .O(new_n4399));
  nor2 g04206(.a(new_n4399), .b(new_n4398), .O(new_n4400));
  nor2 g04207(.a(new_n4400), .b(new_n4289), .O(new_n4401));
  inv1 g04208(.a(new_n4289), .O(new_n4402));
  inv1 g04209(.a(new_n4400), .O(new_n4403));
  nor2 g04210(.a(new_n4403), .b(new_n4402), .O(new_n4404));
  nor2 g04211(.a(new_n4404), .b(new_n4401), .O(new_n4405));
  inv1 g04212(.a(new_n4405), .O(new_n4406));
  nor2 g04213(.a(new_n4406), .b(new_n4200), .O(new_n4407));
  inv1 g04214(.a(new_n4200), .O(new_n4408));
  nor2 g04215(.a(new_n4405), .b(new_n4408), .O(new_n4409));
  nor2 g04216(.a(new_n4409), .b(new_n4407), .O(new_n4410));
  inv1 g04217(.a(new_n4410), .O(new_n4411));
  nor2 g04218(.a(new_n4195), .b(new_n4191), .O(new_n4412));
  nor2 g04219(.a(new_n4412), .b(new_n4411), .O(new_n4413));
  inv1 g04220(.a(new_n4412), .O(new_n4414));
  nor2 g04221(.a(new_n4414), .b(new_n4410), .O(new_n4415));
  nor2 g04222(.a(new_n4415), .b(new_n4413), .O(new_n4416));
  inv1 g04223(.a(new_n4416), .O(\asquared[39] ));
  nor2 g04224(.a(new_n4404), .b(new_n4288), .O(new_n4418));
  nor2 g04225(.a(new_n4398), .b(new_n4323), .O(new_n4419));
  inv1 g04226(.a(new_n4419), .O(new_n4420));
  nor2 g04227(.a(new_n4394), .b(new_n4391), .O(new_n4421));
  nor2 g04228(.a(new_n4314), .b(new_n4309), .O(new_n4422));
  inv1 g04229(.a(new_n4422), .O(new_n4423));
  inv1 g04230(.a(new_n4303), .O(new_n4424));
  inv1 g04231(.a(\a[39] ), .O(new_n4425));
  nor2 g04232(.a(new_n4425), .b(new_n198), .O(new_n4426));
  inv1 g04233(.a(new_n4426), .O(new_n4427));
  nor2 g04234(.a(new_n4427), .b(new_n4424), .O(new_n4428));
  nor2 g04235(.a(new_n4426), .b(new_n4303), .O(new_n4429));
  nor2 g04236(.a(new_n4429), .b(new_n4428), .O(new_n4430));
  inv1 g04237(.a(new_n4430), .O(new_n4431));
  nor2 g04238(.a(new_n1433), .b(new_n4366), .O(new_n4432));
  nor2 g04239(.a(new_n4432), .b(new_n1297), .O(new_n4433));
  nor2 g04240(.a(\a[20] ), .b(new_n194), .O(new_n4434));
  inv1 g04241(.a(new_n4434), .O(new_n4435));
  nor2 g04242(.a(new_n4435), .b(new_n4366), .O(new_n4436));
  nor2 g04243(.a(new_n4436), .b(new_n4433), .O(new_n4437));
  nor2 g04244(.a(new_n4437), .b(new_n4431), .O(new_n4438));
  inv1 g04245(.a(new_n4437), .O(new_n4439));
  nor2 g04246(.a(new_n4439), .b(new_n4430), .O(new_n4440));
  nor2 g04247(.a(new_n4440), .b(new_n4438), .O(new_n4441));
  nor2 g04248(.a(new_n4441), .b(new_n4423), .O(new_n4442));
  inv1 g04249(.a(new_n4441), .O(new_n4443));
  nor2 g04250(.a(new_n4443), .b(new_n4422), .O(new_n4444));
  nor2 g04251(.a(new_n4444), .b(new_n4442), .O(new_n4445));
  nor2 g04252(.a(new_n4214), .b(new_n4208), .O(new_n4446));
  inv1 g04253(.a(new_n4446), .O(new_n4447));
  nor2 g04254(.a(new_n4447), .b(new_n4445), .O(new_n4448));
  inv1 g04255(.a(new_n4445), .O(new_n4449));
  nor2 g04256(.a(new_n4446), .b(new_n4449), .O(new_n4450));
  nor2 g04257(.a(new_n4450), .b(new_n4448), .O(new_n4451));
  inv1 g04258(.a(new_n4451), .O(new_n4452));
  nor2 g04259(.a(new_n4376), .b(new_n4369), .O(new_n4453));
  nor2 g04260(.a(new_n4363), .b(new_n4356), .O(new_n4454));
  nor2 g04261(.a(new_n4454), .b(new_n4453), .O(new_n4455));
  inv1 g04262(.a(new_n4453), .O(new_n4456));
  inv1 g04263(.a(new_n4454), .O(new_n4457));
  nor2 g04264(.a(new_n4457), .b(new_n4456), .O(new_n4458));
  nor2 g04265(.a(new_n4458), .b(new_n4455), .O(new_n4459));
  nor2 g04266(.a(new_n4245), .b(new_n4238), .O(new_n4460));
  nor2 g04267(.a(new_n4460), .b(new_n4459), .O(new_n4461));
  inv1 g04268(.a(new_n4459), .O(new_n4462));
  inv1 g04269(.a(new_n4460), .O(new_n4463));
  nor2 g04270(.a(new_n4463), .b(new_n4462), .O(new_n4464));
  nor2 g04271(.a(new_n4464), .b(new_n4461), .O(new_n4465));
  inv1 g04272(.a(new_n4465), .O(new_n4466));
  nor2 g04273(.a(new_n4266), .b(new_n4260), .O(new_n4467));
  inv1 g04274(.a(new_n4467), .O(new_n4468));
  nor2 g04275(.a(new_n4385), .b(new_n4380), .O(new_n4469));
  inv1 g04276(.a(new_n4469), .O(new_n4470));
  nor2 g04277(.a(new_n4470), .b(new_n4468), .O(new_n4471));
  nor2 g04278(.a(new_n4469), .b(new_n4467), .O(new_n4472));
  nor2 g04279(.a(new_n4472), .b(new_n4471), .O(new_n4473));
  inv1 g04280(.a(new_n4473), .O(new_n4474));
  nor2 g04281(.a(new_n4474), .b(new_n4466), .O(new_n4475));
  nor2 g04282(.a(new_n4473), .b(new_n4465), .O(new_n4476));
  nor2 g04283(.a(new_n4476), .b(new_n4475), .O(new_n4477));
  inv1 g04284(.a(new_n4477), .O(new_n4478));
  nor2 g04285(.a(new_n4478), .b(new_n4452), .O(new_n4479));
  nor2 g04286(.a(new_n4477), .b(new_n4451), .O(new_n4480));
  nor2 g04287(.a(new_n4480), .b(new_n4479), .O(new_n4481));
  inv1 g04288(.a(new_n4481), .O(new_n4482));
  nor2 g04289(.a(new_n4482), .b(new_n4421), .O(new_n4483));
  inv1 g04290(.a(new_n4421), .O(new_n4484));
  nor2 g04291(.a(new_n4481), .b(new_n4484), .O(new_n4485));
  nor2 g04292(.a(new_n4485), .b(new_n4483), .O(new_n4486));
  nor2 g04293(.a(new_n4486), .b(new_n4420), .O(new_n4487));
  inv1 g04294(.a(new_n4486), .O(new_n4488));
  nor2 g04295(.a(new_n4488), .b(new_n4419), .O(new_n4489));
  nor2 g04296(.a(new_n4489), .b(new_n4487), .O(new_n4490));
  inv1 g04297(.a(new_n4490), .O(new_n4491));
  nor2 g04298(.a(new_n4318), .b(new_n4297), .O(new_n4492));
  inv1 g04299(.a(new_n4492), .O(new_n4493));
  nor2 g04300(.a(new_n1736), .b(new_n800), .O(new_n4494));
  nor2 g04301(.a(new_n1647), .b(new_n847), .O(new_n4495));
  nor2 g04302(.a(new_n4495), .b(new_n4494), .O(new_n4496));
  nor2 g04303(.a(new_n1736), .b(new_n847), .O(new_n4497));
  inv1 g04304(.a(new_n4497), .O(new_n4498));
  nor2 g04305(.a(new_n4498), .b(new_n4021), .O(new_n4499));
  nor2 g04306(.a(new_n4499), .b(new_n4496), .O(new_n4500));
  nor2 g04307(.a(new_n4500), .b(new_n4358), .O(new_n4501));
  inv1 g04308(.a(new_n4500), .O(new_n4502));
  nor2 g04309(.a(new_n4502), .b(new_n4357), .O(new_n4503));
  nor2 g04310(.a(new_n4503), .b(new_n4501), .O(new_n4504));
  nor2 g04311(.a(new_n4093), .b(new_n196), .O(new_n4505));
  inv1 g04312(.a(new_n4505), .O(new_n4506));
  nor2 g04313(.a(new_n3870), .b(new_n203), .O(new_n4507));
  nor2 g04314(.a(new_n2121), .b(new_n613), .O(new_n4508));
  nor2 g04315(.a(new_n4508), .b(new_n4507), .O(new_n4509));
  inv1 g04316(.a(new_n4507), .O(new_n4510));
  inv1 g04317(.a(new_n4508), .O(new_n4511));
  nor2 g04318(.a(new_n4511), .b(new_n4510), .O(new_n4512));
  nor2 g04319(.a(new_n4512), .b(new_n4509), .O(new_n4513));
  nor2 g04320(.a(new_n4513), .b(new_n4506), .O(new_n4514));
  inv1 g04321(.a(new_n4513), .O(new_n4515));
  nor2 g04322(.a(new_n4515), .b(new_n4505), .O(new_n4516));
  nor2 g04323(.a(new_n4516), .b(new_n4514), .O(new_n4517));
  nor2 g04324(.a(new_n4517), .b(new_n4504), .O(new_n4518));
  inv1 g04325(.a(new_n4504), .O(new_n4519));
  inv1 g04326(.a(new_n4517), .O(new_n4520));
  nor2 g04327(.a(new_n4520), .b(new_n4519), .O(new_n4521));
  nor2 g04328(.a(new_n4521), .b(new_n4518), .O(new_n4522));
  inv1 g04329(.a(new_n4522), .O(new_n4523));
  nor2 g04330(.a(new_n3231), .b(new_n257), .O(new_n4524));
  inv1 g04331(.a(new_n4524), .O(new_n4525));
  nor2 g04332(.a(new_n2660), .b(new_n363), .O(new_n4526));
  nor2 g04333(.a(new_n3057), .b(new_n295), .O(new_n4527));
  nor2 g04334(.a(new_n4527), .b(new_n4526), .O(new_n4528));
  nor2 g04335(.a(new_n3057), .b(new_n363), .O(new_n4529));
  inv1 g04336(.a(new_n4529), .O(new_n4530));
  nor2 g04337(.a(new_n4530), .b(new_n4227), .O(new_n4531));
  nor2 g04338(.a(new_n4531), .b(new_n4528), .O(new_n4532));
  nor2 g04339(.a(new_n4532), .b(new_n4525), .O(new_n4533));
  inv1 g04340(.a(new_n4532), .O(new_n4534));
  nor2 g04341(.a(new_n4534), .b(new_n4524), .O(new_n4535));
  nor2 g04342(.a(new_n4535), .b(new_n4533), .O(new_n4536));
  nor2 g04343(.a(new_n4536), .b(new_n4523), .O(new_n4537));
  inv1 g04344(.a(new_n4536), .O(new_n4538));
  nor2 g04345(.a(new_n4538), .b(new_n4522), .O(new_n4539));
  nor2 g04346(.a(new_n4539), .b(new_n4537), .O(new_n4540));
  nor2 g04347(.a(new_n4540), .b(new_n4493), .O(new_n4541));
  inv1 g04348(.a(new_n4540), .O(new_n4542));
  nor2 g04349(.a(new_n4542), .b(new_n4492), .O(new_n4543));
  nor2 g04350(.a(new_n4543), .b(new_n4541), .O(new_n4544));
  inv1 g04351(.a(new_n4544), .O(new_n4545));
  nor2 g04352(.a(new_n4271), .b(new_n4220), .O(new_n4546));
  nor2 g04353(.a(new_n4546), .b(new_n4545), .O(new_n4547));
  inv1 g04354(.a(new_n4546), .O(new_n4548));
  nor2 g04355(.a(new_n4548), .b(new_n4544), .O(new_n4549));
  nor2 g04356(.a(new_n4549), .b(new_n4547), .O(new_n4550));
  inv1 g04357(.a(new_n4550), .O(new_n4551));
  nor2 g04358(.a(new_n4283), .b(new_n4277), .O(new_n4552));
  nor2 g04359(.a(new_n4234), .b(new_n4226), .O(new_n4553));
  nor2 g04360(.a(new_n4340), .b(new_n4333), .O(new_n4554));
  nor2 g04361(.a(new_n4554), .b(new_n4553), .O(new_n4555));
  inv1 g04362(.a(new_n4553), .O(new_n4556));
  inv1 g04363(.a(new_n4554), .O(new_n4557));
  nor2 g04364(.a(new_n4557), .b(new_n4556), .O(new_n4558));
  nor2 g04365(.a(new_n4558), .b(new_n4555), .O(new_n4559));
  nor2 g04366(.a(new_n4258), .b(new_n4251), .O(new_n4560));
  nor2 g04367(.a(new_n4560), .b(new_n4559), .O(new_n4561));
  inv1 g04368(.a(new_n4559), .O(new_n4562));
  inv1 g04369(.a(new_n4560), .O(new_n4563));
  nor2 g04370(.a(new_n4563), .b(new_n4562), .O(new_n4564));
  nor2 g04371(.a(new_n4564), .b(new_n4561), .O(new_n4565));
  nor2 g04372(.a(new_n4349), .b(new_n4342), .O(new_n4566));
  inv1 g04373(.a(new_n4566), .O(new_n4567));
  nor2 g04374(.a(new_n4567), .b(new_n4565), .O(new_n4568));
  inv1 g04375(.a(new_n4565), .O(new_n4569));
  nor2 g04376(.a(new_n4566), .b(new_n4569), .O(new_n4570));
  nor2 g04377(.a(new_n4570), .b(new_n4568), .O(new_n4571));
  inv1 g04378(.a(new_n4571), .O(new_n4572));
  nor2 g04379(.a(new_n1297), .b(new_n1199), .O(new_n4573));
  nor2 g04380(.a(new_n1425), .b(new_n1086), .O(new_n4574));
  nor2 g04381(.a(new_n4574), .b(new_n4573), .O(new_n4575));
  nor2 g04382(.a(new_n1425), .b(new_n1199), .O(new_n4576));
  inv1 g04383(.a(new_n4576), .O(new_n4577));
  nor2 g04384(.a(new_n4577), .b(new_n4061), .O(new_n4578));
  nor2 g04385(.a(new_n4578), .b(new_n4575), .O(new_n4579));
  nor2 g04386(.a(new_n4579), .b(new_n4229), .O(new_n4580));
  inv1 g04387(.a(new_n4579), .O(new_n4581));
  nor2 g04388(.a(new_n4581), .b(new_n4228), .O(new_n4582));
  nor2 g04389(.a(new_n4582), .b(new_n4580), .O(new_n4583));
  nor2 g04390(.a(new_n3722), .b(new_n214), .O(new_n4584));
  nor2 g04391(.a(new_n2184), .b(new_n569), .O(new_n4585));
  nor2 g04392(.a(new_n4585), .b(new_n4584), .O(new_n4586));
  inv1 g04393(.a(new_n4584), .O(new_n4587));
  inv1 g04394(.a(new_n4585), .O(new_n4588));
  nor2 g04395(.a(new_n4588), .b(new_n4587), .O(new_n4589));
  nor2 g04396(.a(new_n4589), .b(new_n4586), .O(new_n4590));
  inv1 g04397(.a(new_n4590), .O(new_n4591));
  nor2 g04398(.a(new_n4591), .b(new_n4240), .O(new_n4592));
  nor2 g04399(.a(new_n4590), .b(new_n4239), .O(new_n4593));
  nor2 g04400(.a(new_n4593), .b(new_n4592), .O(new_n4594));
  inv1 g04401(.a(new_n4594), .O(new_n4595));
  nor2 g04402(.a(new_n4595), .b(new_n4583), .O(new_n4596));
  inv1 g04403(.a(new_n4583), .O(new_n4597));
  nor2 g04404(.a(new_n4594), .b(new_n4597), .O(new_n4598));
  nor2 g04405(.a(new_n4598), .b(new_n4596), .O(new_n4599));
  inv1 g04406(.a(new_n4599), .O(new_n4600));
  nor2 g04407(.a(new_n2433), .b(new_n502), .O(new_n4601));
  inv1 g04408(.a(new_n4601), .O(new_n4602));
  nor2 g04409(.a(new_n2506), .b(new_n438), .O(new_n4603));
  nor2 g04410(.a(new_n3533), .b(new_n229), .O(new_n4604));
  nor2 g04411(.a(new_n4604), .b(new_n4603), .O(new_n4605));
  nor2 g04412(.a(new_n3533), .b(new_n438), .O(new_n4606));
  inv1 g04413(.a(new_n4606), .O(new_n4607));
  nor2 g04414(.a(new_n4607), .b(new_n3485), .O(new_n4608));
  nor2 g04415(.a(new_n4608), .b(new_n4605), .O(new_n4609));
  nor2 g04416(.a(new_n4609), .b(new_n4602), .O(new_n4610));
  inv1 g04417(.a(new_n4609), .O(new_n4611));
  nor2 g04418(.a(new_n4611), .b(new_n4601), .O(new_n4612));
  nor2 g04419(.a(new_n4612), .b(new_n4610), .O(new_n4613));
  nor2 g04420(.a(new_n4613), .b(new_n4600), .O(new_n4614));
  inv1 g04421(.a(new_n4613), .O(new_n4615));
  nor2 g04422(.a(new_n4615), .b(new_n4599), .O(new_n4616));
  nor2 g04423(.a(new_n4616), .b(new_n4614), .O(new_n4617));
  inv1 g04424(.a(new_n4617), .O(new_n4618));
  nor2 g04425(.a(new_n4618), .b(new_n4572), .O(new_n4619));
  nor2 g04426(.a(new_n4617), .b(new_n4571), .O(new_n4620));
  nor2 g04427(.a(new_n4620), .b(new_n4619), .O(new_n4621));
  inv1 g04428(.a(new_n4621), .O(new_n4622));
  nor2 g04429(.a(new_n4622), .b(new_n4552), .O(new_n4623));
  inv1 g04430(.a(new_n4552), .O(new_n4624));
  nor2 g04431(.a(new_n4621), .b(new_n4624), .O(new_n4625));
  nor2 g04432(.a(new_n4625), .b(new_n4623), .O(new_n4626));
  inv1 g04433(.a(new_n4626), .O(new_n4627));
  nor2 g04434(.a(new_n4627), .b(new_n4551), .O(new_n4628));
  nor2 g04435(.a(new_n4626), .b(new_n4550), .O(new_n4629));
  nor2 g04436(.a(new_n4629), .b(new_n4628), .O(new_n4630));
  inv1 g04437(.a(new_n4630), .O(new_n4631));
  nor2 g04438(.a(new_n4631), .b(new_n4491), .O(new_n4632));
  nor2 g04439(.a(new_n4630), .b(new_n4490), .O(new_n4633));
  nor2 g04440(.a(new_n4633), .b(new_n4632), .O(new_n4634));
  inv1 g04441(.a(new_n4634), .O(new_n4635));
  nor2 g04442(.a(new_n4635), .b(new_n4418), .O(new_n4636));
  inv1 g04443(.a(new_n4418), .O(new_n4637));
  nor2 g04444(.a(new_n4634), .b(new_n4637), .O(new_n4638));
  nor2 g04445(.a(new_n4638), .b(new_n4636), .O(new_n4639));
  inv1 g04446(.a(new_n4639), .O(new_n4640));
  nor2 g04447(.a(new_n4413), .b(new_n4409), .O(new_n4641));
  nor2 g04448(.a(new_n4641), .b(new_n4640), .O(new_n4642));
  inv1 g04449(.a(new_n4641), .O(new_n4643));
  nor2 g04450(.a(new_n4643), .b(new_n4639), .O(new_n4644));
  nor2 g04451(.a(new_n4644), .b(new_n4642), .O(new_n4645));
  inv1 g04452(.a(new_n4645), .O(\asquared[40] ));
  nor2 g04453(.a(new_n4632), .b(new_n4489), .O(new_n4647));
  nor2 g04454(.a(new_n4503), .b(new_n4496), .O(new_n4648));
  nor2 g04455(.a(new_n4535), .b(new_n4528), .O(new_n4649));
  nor2 g04456(.a(new_n4649), .b(new_n4648), .O(new_n4650));
  inv1 g04457(.a(new_n4648), .O(new_n4651));
  inv1 g04458(.a(new_n4649), .O(new_n4652));
  nor2 g04459(.a(new_n4652), .b(new_n4651), .O(new_n4653));
  nor2 g04460(.a(new_n4653), .b(new_n4650), .O(new_n4654));
  nor2 g04461(.a(new_n4438), .b(new_n4428), .O(new_n4655));
  inv1 g04462(.a(new_n4655), .O(new_n4656));
  nor2 g04463(.a(new_n4656), .b(new_n4654), .O(new_n4657));
  inv1 g04464(.a(new_n4654), .O(new_n4658));
  nor2 g04465(.a(new_n4655), .b(new_n4658), .O(new_n4659));
  nor2 g04466(.a(new_n4659), .b(new_n4657), .O(new_n4660));
  nor2 g04467(.a(new_n4450), .b(new_n4444), .O(new_n4661));
  inv1 g04468(.a(new_n4661), .O(new_n4662));
  nor2 g04469(.a(new_n4662), .b(new_n4660), .O(new_n4663));
  inv1 g04470(.a(new_n4660), .O(new_n4664));
  nor2 g04471(.a(new_n4661), .b(new_n4664), .O(new_n4665));
  nor2 g04472(.a(new_n4665), .b(new_n4663), .O(new_n4666));
  nor2 g04473(.a(new_n3870), .b(new_n214), .O(new_n4667));
  inv1 g04474(.a(new_n4667), .O(new_n4668));
  nor2 g04475(.a(new_n2433), .b(new_n569), .O(new_n4669));
  nor2 g04476(.a(new_n3722), .b(new_n229), .O(new_n4670));
  nor2 g04477(.a(new_n4670), .b(new_n4669), .O(new_n4671));
  inv1 g04478(.a(new_n4669), .O(new_n4672));
  inv1 g04479(.a(new_n4670), .O(new_n4673));
  nor2 g04480(.a(new_n4673), .b(new_n4672), .O(new_n4674));
  nor2 g04481(.a(new_n4674), .b(new_n4671), .O(new_n4675));
  nor2 g04482(.a(new_n4675), .b(new_n4668), .O(new_n4676));
  inv1 g04483(.a(new_n4675), .O(new_n4677));
  nor2 g04484(.a(new_n4677), .b(new_n4667), .O(new_n4678));
  nor2 g04485(.a(new_n4678), .b(new_n4676), .O(new_n4679));
  inv1 g04486(.a(new_n4679), .O(new_n4680));
  nor2 g04487(.a(new_n1493), .b(new_n1086), .O(new_n4681));
  inv1 g04488(.a(\a[40] ), .O(new_n4682));
  nor2 g04489(.a(new_n4682), .b(new_n198), .O(new_n4683));
  nor2 g04490(.a(new_n4683), .b(new_n4370), .O(new_n4684));
  inv1 g04491(.a(new_n4367), .O(new_n4685));
  nor2 g04492(.a(new_n4682), .b(new_n196), .O(new_n4686));
  inv1 g04493(.a(new_n4686), .O(new_n4687));
  nor2 g04494(.a(new_n4687), .b(new_n4685), .O(new_n4688));
  nor2 g04495(.a(new_n4688), .b(new_n4684), .O(new_n4689));
  inv1 g04496(.a(new_n4689), .O(new_n4690));
  nor2 g04497(.a(new_n4690), .b(new_n4681), .O(new_n4691));
  inv1 g04498(.a(new_n4681), .O(new_n4692));
  nor2 g04499(.a(new_n4689), .b(new_n4692), .O(new_n4693));
  nor2 g04500(.a(new_n4693), .b(new_n4691), .O(new_n4694));
  nor2 g04501(.a(new_n3231), .b(new_n295), .O(new_n4695));
  inv1 g04502(.a(new_n4695), .O(new_n4696));
  nor2 g04503(.a(new_n3057), .b(new_n322), .O(new_n4697));
  nor2 g04504(.a(new_n4697), .b(new_n2830), .O(new_n4698));
  nor2 g04505(.a(new_n4530), .b(new_n4229), .O(new_n4699));
  nor2 g04506(.a(new_n4699), .b(new_n4698), .O(new_n4700));
  nor2 g04507(.a(new_n4700), .b(new_n4696), .O(new_n4701));
  inv1 g04508(.a(new_n4700), .O(new_n4702));
  nor2 g04509(.a(new_n4702), .b(new_n4695), .O(new_n4703));
  nor2 g04510(.a(new_n4703), .b(new_n4701), .O(new_n4704));
  nor2 g04511(.a(new_n4704), .b(new_n4694), .O(new_n4705));
  inv1 g04512(.a(new_n4694), .O(new_n4706));
  inv1 g04513(.a(new_n4704), .O(new_n4707));
  nor2 g04514(.a(new_n4707), .b(new_n4706), .O(new_n4708));
  nor2 g04515(.a(new_n4708), .b(new_n4705), .O(new_n4709));
  nor2 g04516(.a(new_n4709), .b(new_n4680), .O(new_n4710));
  inv1 g04517(.a(new_n4709), .O(new_n4711));
  nor2 g04518(.a(new_n4711), .b(new_n4679), .O(new_n4712));
  nor2 g04519(.a(new_n4712), .b(new_n4710), .O(new_n4713));
  nor2 g04520(.a(new_n4713), .b(new_n4666), .O(new_n4714));
  inv1 g04521(.a(new_n4666), .O(new_n4715));
  inv1 g04522(.a(new_n4713), .O(new_n4716));
  nor2 g04523(.a(new_n4716), .b(new_n4715), .O(new_n4717));
  nor2 g04524(.a(new_n4717), .b(new_n4714), .O(new_n4718));
  inv1 g04525(.a(new_n4718), .O(new_n4719));
  nor2 g04526(.a(new_n4483), .b(new_n4479), .O(new_n4720));
  nor2 g04527(.a(new_n4720), .b(new_n4719), .O(new_n4721));
  inv1 g04528(.a(new_n4720), .O(new_n4722));
  nor2 g04529(.a(new_n4722), .b(new_n4718), .O(new_n4723));
  nor2 g04530(.a(new_n4723), .b(new_n4721), .O(new_n4724));
  inv1 g04531(.a(new_n4724), .O(new_n4725));
  nor2 g04532(.a(new_n4475), .b(new_n4472), .O(new_n4726));
  nor2 g04533(.a(new_n2506), .b(new_n502), .O(new_n4727));
  inv1 g04534(.a(new_n4727), .O(new_n4728));
  nor2 g04535(.a(new_n3533), .b(new_n257), .O(new_n4729));
  nor2 g04536(.a(new_n2660), .b(new_n438), .O(new_n4730));
  nor2 g04537(.a(new_n4730), .b(new_n4729), .O(new_n4731));
  inv1 g04538(.a(new_n4729), .O(new_n4732));
  inv1 g04539(.a(new_n4730), .O(new_n4733));
  nor2 g04540(.a(new_n4733), .b(new_n4732), .O(new_n4734));
  nor2 g04541(.a(new_n4734), .b(new_n4731), .O(new_n4735));
  nor2 g04542(.a(new_n4735), .b(new_n4728), .O(new_n4736));
  inv1 g04543(.a(new_n4735), .O(new_n4737));
  nor2 g04544(.a(new_n4737), .b(new_n4727), .O(new_n4738));
  nor2 g04545(.a(new_n4738), .b(new_n4736), .O(new_n4739));
  inv1 g04546(.a(new_n4739), .O(new_n4740));
  nor2 g04547(.a(new_n4093), .b(new_n203), .O(new_n4741));
  nor2 g04548(.a(new_n2184), .b(new_n613), .O(new_n4742));
  nor2 g04549(.a(new_n2121), .b(new_n699), .O(new_n4743));
  nor2 g04550(.a(new_n4743), .b(new_n4742), .O(new_n4744));
  nor2 g04551(.a(new_n2184), .b(new_n699), .O(new_n4745));
  inv1 g04552(.a(new_n4745), .O(new_n4746));
  nor2 g04553(.a(new_n4746), .b(new_n4511), .O(new_n4747));
  nor2 g04554(.a(new_n4747), .b(new_n4744), .O(new_n4748));
  inv1 g04555(.a(new_n4748), .O(new_n4749));
  nor2 g04556(.a(new_n4749), .b(new_n4741), .O(new_n4750));
  inv1 g04557(.a(new_n4741), .O(new_n4751));
  nor2 g04558(.a(new_n4748), .b(new_n4751), .O(new_n4752));
  nor2 g04559(.a(new_n4752), .b(new_n4750), .O(new_n4753));
  nor2 g04560(.a(new_n1903), .b(new_n800), .O(new_n4754));
  inv1 g04561(.a(new_n4754), .O(new_n4755));
  nor2 g04562(.a(new_n1647), .b(new_n941), .O(new_n4756));
  nor2 g04563(.a(new_n4756), .b(new_n4497), .O(new_n4757));
  inv1 g04564(.a(new_n4495), .O(new_n4758));
  nor2 g04565(.a(new_n1736), .b(new_n941), .O(new_n4759));
  inv1 g04566(.a(new_n4759), .O(new_n4760));
  nor2 g04567(.a(new_n4760), .b(new_n4758), .O(new_n4761));
  nor2 g04568(.a(new_n4761), .b(new_n4757), .O(new_n4762));
  nor2 g04569(.a(new_n4762), .b(new_n4755), .O(new_n4763));
  inv1 g04570(.a(new_n4762), .O(new_n4764));
  nor2 g04571(.a(new_n4764), .b(new_n4754), .O(new_n4765));
  nor2 g04572(.a(new_n4765), .b(new_n4763), .O(new_n4766));
  nor2 g04573(.a(new_n4766), .b(new_n4753), .O(new_n4767));
  inv1 g04574(.a(new_n4753), .O(new_n4768));
  inv1 g04575(.a(new_n4766), .O(new_n4769));
  nor2 g04576(.a(new_n4769), .b(new_n4768), .O(new_n4770));
  nor2 g04577(.a(new_n4770), .b(new_n4767), .O(new_n4771));
  nor2 g04578(.a(new_n4771), .b(new_n4740), .O(new_n4772));
  inv1 g04579(.a(new_n4771), .O(new_n4773));
  nor2 g04580(.a(new_n4773), .b(new_n4739), .O(new_n4774));
  nor2 g04581(.a(new_n4774), .b(new_n4772), .O(new_n4775));
  inv1 g04582(.a(new_n4775), .O(new_n4776));
  nor2 g04583(.a(new_n4776), .b(new_n4726), .O(new_n4777));
  inv1 g04584(.a(new_n4726), .O(new_n4778));
  nor2 g04585(.a(new_n4775), .b(new_n4778), .O(new_n4779));
  nor2 g04586(.a(new_n4779), .b(new_n4777), .O(new_n4780));
  inv1 g04587(.a(new_n4780), .O(new_n4781));
  nor2 g04588(.a(new_n4564), .b(new_n4558), .O(new_n4782));
  inv1 g04589(.a(new_n4782), .O(new_n4783));
  nor2 g04590(.a(new_n4464), .b(new_n4458), .O(new_n4784));
  inv1 g04591(.a(new_n4784), .O(new_n4785));
  nor2 g04592(.a(new_n4785), .b(new_n4783), .O(new_n4786));
  nor2 g04593(.a(new_n4784), .b(new_n4782), .O(new_n4787));
  nor2 g04594(.a(new_n4787), .b(new_n4786), .O(new_n4788));
  inv1 g04595(.a(new_n4788), .O(new_n4789));
  inv1 g04596(.a(new_n4432), .O(new_n4790));
  nor2 g04597(.a(new_n4425), .b(new_n194), .O(new_n4791));
  nor2 g04598(.a(new_n4791), .b(new_n4576), .O(new_n4792));
  inv1 g04599(.a(new_n4791), .O(new_n4793));
  nor2 g04600(.a(new_n4793), .b(new_n4577), .O(new_n4794));
  nor2 g04601(.a(new_n4794), .b(new_n4792), .O(new_n4795));
  inv1 g04602(.a(new_n4795), .O(new_n4796));
  nor2 g04603(.a(new_n4796), .b(new_n4790), .O(new_n4797));
  nor2 g04604(.a(new_n4795), .b(new_n4432), .O(new_n4798));
  nor2 g04605(.a(new_n4798), .b(new_n4797), .O(new_n4799));
  inv1 g04606(.a(new_n4799), .O(new_n4800));
  nor2 g04607(.a(new_n4582), .b(new_n4575), .O(new_n4801));
  inv1 g04608(.a(new_n4801), .O(new_n4802));
  nor2 g04609(.a(new_n4802), .b(new_n4800), .O(new_n4803));
  nor2 g04610(.a(new_n4801), .b(new_n4799), .O(new_n4804));
  nor2 g04611(.a(new_n4804), .b(new_n4803), .O(new_n4805));
  inv1 g04612(.a(new_n4805), .O(new_n4806));
  nor2 g04613(.a(new_n4806), .b(new_n4789), .O(new_n4807));
  nor2 g04614(.a(new_n4805), .b(new_n4788), .O(new_n4808));
  nor2 g04615(.a(new_n4808), .b(new_n4807), .O(new_n4809));
  inv1 g04616(.a(new_n4809), .O(new_n4810));
  nor2 g04617(.a(new_n4810), .b(new_n4781), .O(new_n4811));
  nor2 g04618(.a(new_n4809), .b(new_n4780), .O(new_n4812));
  nor2 g04619(.a(new_n4812), .b(new_n4811), .O(new_n4813));
  inv1 g04620(.a(new_n4813), .O(new_n4814));
  nor2 g04621(.a(new_n4814), .b(new_n4725), .O(new_n4815));
  nor2 g04622(.a(new_n4813), .b(new_n4724), .O(new_n4816));
  nor2 g04623(.a(new_n4816), .b(new_n4815), .O(new_n4817));
  inv1 g04624(.a(new_n4817), .O(new_n4818));
  nor2 g04625(.a(new_n4547), .b(new_n4543), .O(new_n4819));
  nor2 g04626(.a(new_n4619), .b(new_n4570), .O(new_n4820));
  nor2 g04627(.a(new_n4592), .b(new_n4589), .O(new_n4821));
  inv1 g04628(.a(new_n4821), .O(new_n4822));
  nor2 g04629(.a(new_n4516), .b(new_n4509), .O(new_n4823));
  nor2 g04630(.a(new_n4612), .b(new_n4605), .O(new_n4824));
  nor2 g04631(.a(new_n4824), .b(new_n4823), .O(new_n4825));
  inv1 g04632(.a(new_n4823), .O(new_n4826));
  inv1 g04633(.a(new_n4824), .O(new_n4827));
  nor2 g04634(.a(new_n4827), .b(new_n4826), .O(new_n4828));
  nor2 g04635(.a(new_n4828), .b(new_n4825), .O(new_n4829));
  nor2 g04636(.a(new_n4829), .b(new_n4822), .O(new_n4830));
  inv1 g04637(.a(new_n4829), .O(new_n4831));
  nor2 g04638(.a(new_n4831), .b(new_n4821), .O(new_n4832));
  nor2 g04639(.a(new_n4832), .b(new_n4830), .O(new_n4833));
  inv1 g04640(.a(new_n4833), .O(new_n4834));
  nor2 g04641(.a(new_n4614), .b(new_n4596), .O(new_n4835));
  inv1 g04642(.a(new_n4835), .O(new_n4836));
  nor2 g04643(.a(new_n4537), .b(new_n4518), .O(new_n4837));
  inv1 g04644(.a(new_n4837), .O(new_n4838));
  nor2 g04645(.a(new_n4838), .b(new_n4836), .O(new_n4839));
  nor2 g04646(.a(new_n4837), .b(new_n4835), .O(new_n4840));
  nor2 g04647(.a(new_n4840), .b(new_n4839), .O(new_n4841));
  inv1 g04648(.a(new_n4841), .O(new_n4842));
  nor2 g04649(.a(new_n4842), .b(new_n4834), .O(new_n4843));
  nor2 g04650(.a(new_n4841), .b(new_n4833), .O(new_n4844));
  nor2 g04651(.a(new_n4844), .b(new_n4843), .O(new_n4845));
  inv1 g04652(.a(new_n4845), .O(new_n4846));
  nor2 g04653(.a(new_n4846), .b(new_n4820), .O(new_n4847));
  inv1 g04654(.a(new_n4820), .O(new_n4848));
  nor2 g04655(.a(new_n4845), .b(new_n4848), .O(new_n4849));
  nor2 g04656(.a(new_n4849), .b(new_n4847), .O(new_n4850));
  inv1 g04657(.a(new_n4850), .O(new_n4851));
  nor2 g04658(.a(new_n4851), .b(new_n4819), .O(new_n4852));
  inv1 g04659(.a(new_n4819), .O(new_n4853));
  nor2 g04660(.a(new_n4850), .b(new_n4853), .O(new_n4854));
  nor2 g04661(.a(new_n4854), .b(new_n4852), .O(new_n4855));
  inv1 g04662(.a(new_n4855), .O(new_n4856));
  nor2 g04663(.a(new_n4628), .b(new_n4623), .O(new_n4857));
  nor2 g04664(.a(new_n4857), .b(new_n4856), .O(new_n4858));
  inv1 g04665(.a(new_n4857), .O(new_n4859));
  nor2 g04666(.a(new_n4859), .b(new_n4855), .O(new_n4860));
  nor2 g04667(.a(new_n4860), .b(new_n4858), .O(new_n4861));
  inv1 g04668(.a(new_n4861), .O(new_n4862));
  nor2 g04669(.a(new_n4862), .b(new_n4818), .O(new_n4863));
  nor2 g04670(.a(new_n4861), .b(new_n4817), .O(new_n4864));
  nor2 g04671(.a(new_n4864), .b(new_n4863), .O(new_n4865));
  inv1 g04672(.a(new_n4865), .O(new_n4866));
  nor2 g04673(.a(new_n4866), .b(new_n4647), .O(new_n4867));
  inv1 g04674(.a(new_n4647), .O(new_n4868));
  nor2 g04675(.a(new_n4865), .b(new_n4868), .O(new_n4869));
  nor2 g04676(.a(new_n4869), .b(new_n4867), .O(new_n4870));
  inv1 g04677(.a(new_n4870), .O(new_n4871));
  nor2 g04678(.a(new_n4642), .b(new_n4638), .O(new_n4872));
  nor2 g04679(.a(new_n4872), .b(new_n4871), .O(new_n4873));
  inv1 g04680(.a(new_n4872), .O(new_n4874));
  nor2 g04681(.a(new_n4874), .b(new_n4870), .O(new_n4875));
  nor2 g04682(.a(new_n4875), .b(new_n4873), .O(new_n4876));
  inv1 g04683(.a(new_n4876), .O(\asquared[41] ));
  nor2 g04684(.a(new_n4863), .b(new_n4858), .O(new_n4878));
  inv1 g04685(.a(new_n4878), .O(new_n4879));
  nor2 g04686(.a(new_n4811), .b(new_n4777), .O(new_n4880));
  inv1 g04687(.a(new_n4880), .O(new_n4881));
  nor2 g04688(.a(new_n4717), .b(new_n4665), .O(new_n4882));
  nor2 g04689(.a(new_n4765), .b(new_n4757), .O(new_n4883));
  nor2 g04690(.a(new_n4691), .b(new_n4684), .O(new_n4884));
  nor2 g04691(.a(new_n4884), .b(new_n4883), .O(new_n4885));
  inv1 g04692(.a(new_n4883), .O(new_n4886));
  inv1 g04693(.a(new_n4884), .O(new_n4887));
  nor2 g04694(.a(new_n4887), .b(new_n4886), .O(new_n4888));
  nor2 g04695(.a(new_n4888), .b(new_n4885), .O(new_n4889));
  nor2 g04696(.a(new_n4750), .b(new_n4744), .O(new_n4890));
  nor2 g04697(.a(new_n4890), .b(new_n4889), .O(new_n4891));
  inv1 g04698(.a(new_n4889), .O(new_n4892));
  inv1 g04699(.a(new_n4890), .O(new_n4893));
  nor2 g04700(.a(new_n4893), .b(new_n4892), .O(new_n4894));
  nor2 g04701(.a(new_n4894), .b(new_n4891), .O(new_n4895));
  nor2 g04702(.a(new_n4712), .b(new_n4705), .O(new_n4896));
  inv1 g04703(.a(new_n4896), .O(new_n4897));
  nor2 g04704(.a(new_n4897), .b(new_n4895), .O(new_n4898));
  inv1 g04705(.a(new_n4895), .O(new_n4899));
  nor2 g04706(.a(new_n4896), .b(new_n4899), .O(new_n4900));
  nor2 g04707(.a(new_n4900), .b(new_n4898), .O(new_n4901));
  inv1 g04708(.a(new_n4901), .O(new_n4902));
  nor2 g04709(.a(new_n1550), .b(new_n4682), .O(new_n4903));
  nor2 g04710(.a(new_n4682), .b(new_n194), .O(new_n4904));
  nor2 g04711(.a(new_n4904), .b(\a[21] ), .O(new_n4905));
  nor2 g04712(.a(new_n4905), .b(new_n4903), .O(new_n4906));
  nor2 g04713(.a(new_n4703), .b(new_n4698), .O(new_n4907));
  nor2 g04714(.a(new_n4907), .b(new_n4906), .O(new_n4908));
  inv1 g04715(.a(new_n4906), .O(new_n4909));
  inv1 g04716(.a(new_n4907), .O(new_n4910));
  nor2 g04717(.a(new_n4910), .b(new_n4909), .O(new_n4911));
  nor2 g04718(.a(new_n4911), .b(new_n4908), .O(new_n4912));
  inv1 g04719(.a(new_n4912), .O(new_n4913));
  nor2 g04720(.a(new_n4738), .b(new_n4731), .O(new_n4914));
  inv1 g04721(.a(new_n4914), .O(new_n4915));
  nor2 g04722(.a(new_n4915), .b(new_n4913), .O(new_n4916));
  nor2 g04723(.a(new_n4914), .b(new_n4912), .O(new_n4917));
  nor2 g04724(.a(new_n4917), .b(new_n4916), .O(new_n4918));
  inv1 g04725(.a(new_n4918), .O(new_n4919));
  nor2 g04726(.a(new_n4919), .b(new_n4902), .O(new_n4920));
  nor2 g04727(.a(new_n4918), .b(new_n4901), .O(new_n4921));
  nor2 g04728(.a(new_n4921), .b(new_n4920), .O(new_n4922));
  inv1 g04729(.a(new_n4922), .O(new_n4923));
  nor2 g04730(.a(new_n4923), .b(new_n4882), .O(new_n4924));
  inv1 g04731(.a(new_n4882), .O(new_n4925));
  nor2 g04732(.a(new_n4922), .b(new_n4925), .O(new_n4926));
  nor2 g04733(.a(new_n4926), .b(new_n4924), .O(new_n4927));
  nor2 g04734(.a(new_n4927), .b(new_n4881), .O(new_n4928));
  inv1 g04735(.a(new_n4927), .O(new_n4929));
  nor2 g04736(.a(new_n4929), .b(new_n4880), .O(new_n4930));
  nor2 g04737(.a(new_n4930), .b(new_n4928), .O(new_n4931));
  nor2 g04738(.a(new_n4815), .b(new_n4721), .O(new_n4932));
  inv1 g04739(.a(new_n4932), .O(new_n4933));
  nor2 g04740(.a(new_n4933), .b(new_n4931), .O(new_n4934));
  inv1 g04741(.a(new_n4931), .O(new_n4935));
  nor2 g04742(.a(new_n4932), .b(new_n4935), .O(new_n4936));
  nor2 g04743(.a(new_n4936), .b(new_n4934), .O(new_n4937));
  inv1 g04744(.a(new_n4937), .O(new_n4938));
  nor2 g04745(.a(new_n4659), .b(new_n4653), .O(new_n4939));
  inv1 g04746(.a(new_n4939), .O(new_n4940));
  nor2 g04747(.a(new_n4832), .b(new_n4828), .O(new_n4941));
  inv1 g04748(.a(new_n4941), .O(new_n4942));
  nor2 g04749(.a(new_n4942), .b(new_n4940), .O(new_n4943));
  nor2 g04750(.a(new_n4941), .b(new_n4939), .O(new_n4944));
  nor2 g04751(.a(new_n4944), .b(new_n4943), .O(new_n4945));
  nor2 g04752(.a(new_n4774), .b(new_n4767), .O(new_n4946));
  inv1 g04753(.a(new_n4946), .O(new_n4947));
  nor2 g04754(.a(new_n4947), .b(new_n4945), .O(new_n4948));
  inv1 g04755(.a(new_n4945), .O(new_n4949));
  nor2 g04756(.a(new_n4946), .b(new_n4949), .O(new_n4950));
  nor2 g04757(.a(new_n4950), .b(new_n4948), .O(new_n4951));
  nor2 g04758(.a(new_n4843), .b(new_n4840), .O(new_n4952));
  inv1 g04759(.a(new_n4794), .O(new_n4953));
  inv1 g04760(.a(\a[41] ), .O(new_n4954));
  nor2 g04761(.a(new_n4954), .b(new_n198), .O(new_n4955));
  nor2 g04762(.a(new_n4425), .b(new_n196), .O(new_n4956));
  nor2 g04763(.a(new_n4956), .b(new_n4955), .O(new_n4957));
  nor2 g04764(.a(new_n4954), .b(new_n196), .O(new_n4958));
  inv1 g04765(.a(new_n4958), .O(new_n4959));
  nor2 g04766(.a(new_n4959), .b(new_n4427), .O(new_n4960));
  nor2 g04767(.a(new_n4960), .b(new_n4957), .O(new_n4961));
  inv1 g04768(.a(new_n4961), .O(new_n4962));
  nor2 g04769(.a(new_n4962), .b(new_n4953), .O(new_n4963));
  nor2 g04770(.a(new_n4961), .b(new_n4794), .O(new_n4964));
  nor2 g04771(.a(new_n4964), .b(new_n4963), .O(new_n4965));
  inv1 g04772(.a(new_n4965), .O(new_n4966));
  nor2 g04773(.a(new_n4678), .b(new_n4671), .O(new_n4967));
  inv1 g04774(.a(new_n4967), .O(new_n4968));
  nor2 g04775(.a(new_n4968), .b(new_n4966), .O(new_n4969));
  nor2 g04776(.a(new_n4967), .b(new_n4965), .O(new_n4970));
  nor2 g04777(.a(new_n4970), .b(new_n4969), .O(new_n4971));
  inv1 g04778(.a(new_n4971), .O(new_n4972));
  nor2 g04779(.a(new_n4366), .b(new_n203), .O(new_n4973));
  inv1 g04780(.a(new_n4973), .O(new_n4974));
  nor2 g04781(.a(new_n2433), .b(new_n613), .O(new_n4975));
  nor2 g04782(.a(new_n2121), .b(new_n800), .O(new_n4976));
  nor2 g04783(.a(new_n4976), .b(new_n4975), .O(new_n4977));
  nor2 g04784(.a(new_n2433), .b(new_n800), .O(new_n4978));
  inv1 g04785(.a(new_n4978), .O(new_n4979));
  nor2 g04786(.a(new_n4979), .b(new_n4511), .O(new_n4980));
  nor2 g04787(.a(new_n4980), .b(new_n4977), .O(new_n4981));
  nor2 g04788(.a(new_n4981), .b(new_n4974), .O(new_n4982));
  inv1 g04789(.a(new_n4981), .O(new_n4983));
  nor2 g04790(.a(new_n4983), .b(new_n4973), .O(new_n4984));
  nor2 g04791(.a(new_n4984), .b(new_n4982), .O(new_n4985));
  nor2 g04792(.a(new_n4985), .b(new_n4972), .O(new_n4986));
  inv1 g04793(.a(new_n4985), .O(new_n4987));
  nor2 g04794(.a(new_n4987), .b(new_n4971), .O(new_n4988));
  nor2 g04795(.a(new_n4988), .b(new_n4986), .O(new_n4989));
  inv1 g04796(.a(new_n4989), .O(new_n4990));
  nor2 g04797(.a(new_n4990), .b(new_n4952), .O(new_n4991));
  inv1 g04798(.a(new_n4952), .O(new_n4992));
  nor2 g04799(.a(new_n4989), .b(new_n4992), .O(new_n4993));
  nor2 g04800(.a(new_n4993), .b(new_n4991), .O(new_n4994));
  nor2 g04801(.a(new_n4994), .b(new_n4951), .O(new_n4995));
  inv1 g04802(.a(new_n4951), .O(new_n4996));
  inv1 g04803(.a(new_n4994), .O(new_n4997));
  nor2 g04804(.a(new_n4997), .b(new_n4996), .O(new_n4998));
  nor2 g04805(.a(new_n4998), .b(new_n4995), .O(new_n4999));
  inv1 g04806(.a(new_n4999), .O(new_n5000));
  nor2 g04807(.a(new_n4852), .b(new_n4847), .O(new_n5001));
  nor2 g04808(.a(new_n4803), .b(new_n4797), .O(new_n5002));
  inv1 g04809(.a(new_n5002), .O(new_n5003));
  nor2 g04810(.a(new_n3870), .b(new_n229), .O(new_n5004));
  nor2 g04811(.a(new_n3722), .b(new_n257), .O(new_n5005));
  nor2 g04812(.a(new_n2660), .b(new_n502), .O(new_n5006));
  nor2 g04813(.a(new_n5006), .b(new_n5005), .O(new_n5007));
  nor2 g04814(.a(new_n3722), .b(new_n502), .O(new_n5008));
  inv1 g04815(.a(new_n5008), .O(new_n5009));
  nor2 g04816(.a(new_n5009), .b(new_n3922), .O(new_n5010));
  nor2 g04817(.a(new_n5010), .b(new_n5007), .O(new_n5011));
  inv1 g04818(.a(new_n5011), .O(new_n5012));
  nor2 g04819(.a(new_n5012), .b(new_n5004), .O(new_n5013));
  inv1 g04820(.a(new_n5004), .O(new_n5014));
  nor2 g04821(.a(new_n5011), .b(new_n5014), .O(new_n5015));
  nor2 g04822(.a(new_n5015), .b(new_n5013), .O(new_n5016));
  nor2 g04823(.a(new_n3231), .b(new_n322), .O(new_n5017));
  inv1 g04824(.a(new_n5017), .O(new_n5018));
  nor2 g04825(.a(new_n1425), .b(new_n1297), .O(new_n5019));
  nor2 g04826(.a(new_n1493), .b(new_n1199), .O(new_n5020));
  nor2 g04827(.a(new_n5020), .b(new_n5019), .O(new_n5021));
  inv1 g04828(.a(new_n5019), .O(new_n5022));
  inv1 g04829(.a(new_n5020), .O(new_n5023));
  nor2 g04830(.a(new_n5023), .b(new_n5022), .O(new_n5024));
  nor2 g04831(.a(new_n5024), .b(new_n5021), .O(new_n5025));
  nor2 g04832(.a(new_n5025), .b(new_n5018), .O(new_n5026));
  inv1 g04833(.a(new_n5025), .O(new_n5027));
  nor2 g04834(.a(new_n5027), .b(new_n5017), .O(new_n5028));
  nor2 g04835(.a(new_n5028), .b(new_n5026), .O(new_n5029));
  nor2 g04836(.a(new_n5029), .b(new_n5016), .O(new_n5030));
  inv1 g04837(.a(new_n5016), .O(new_n5031));
  inv1 g04838(.a(new_n5029), .O(new_n5032));
  nor2 g04839(.a(new_n5032), .b(new_n5031), .O(new_n5033));
  nor2 g04840(.a(new_n5033), .b(new_n5030), .O(new_n5034));
  nor2 g04841(.a(new_n5034), .b(new_n5003), .O(new_n5035));
  inv1 g04842(.a(new_n5034), .O(new_n5036));
  nor2 g04843(.a(new_n5036), .b(new_n5002), .O(new_n5037));
  nor2 g04844(.a(new_n5037), .b(new_n5035), .O(new_n5038));
  nor2 g04845(.a(new_n4807), .b(new_n4787), .O(new_n5039));
  inv1 g04846(.a(new_n5039), .O(new_n5040));
  nor2 g04847(.a(new_n5040), .b(new_n5038), .O(new_n5041));
  inv1 g04848(.a(new_n5038), .O(new_n5042));
  nor2 g04849(.a(new_n5039), .b(new_n5042), .O(new_n5043));
  nor2 g04850(.a(new_n5043), .b(new_n5041), .O(new_n5044));
  nor2 g04851(.a(new_n1903), .b(new_n847), .O(new_n5045));
  inv1 g04852(.a(new_n5045), .O(new_n5046));
  nor2 g04853(.a(new_n1647), .b(new_n1086), .O(new_n5047));
  nor2 g04854(.a(new_n5047), .b(new_n4759), .O(new_n5048));
  inv1 g04855(.a(new_n4756), .O(new_n5049));
  nor2 g04856(.a(new_n1736), .b(new_n1086), .O(new_n5050));
  inv1 g04857(.a(new_n5050), .O(new_n5051));
  nor2 g04858(.a(new_n5051), .b(new_n5049), .O(new_n5052));
  nor2 g04859(.a(new_n5052), .b(new_n5048), .O(new_n5053));
  nor2 g04860(.a(new_n5053), .b(new_n5046), .O(new_n5054));
  inv1 g04861(.a(new_n5053), .O(new_n5055));
  nor2 g04862(.a(new_n5055), .b(new_n5045), .O(new_n5056));
  nor2 g04863(.a(new_n5056), .b(new_n5054), .O(new_n5057));
  nor2 g04864(.a(new_n4093), .b(new_n214), .O(new_n5058));
  nor2 g04865(.a(new_n2506), .b(new_n569), .O(new_n5059));
  nor2 g04866(.a(new_n5059), .b(new_n5058), .O(new_n5060));
  inv1 g04867(.a(new_n5058), .O(new_n5061));
  inv1 g04868(.a(new_n5059), .O(new_n5062));
  nor2 g04869(.a(new_n5062), .b(new_n5061), .O(new_n5063));
  nor2 g04870(.a(new_n5063), .b(new_n5060), .O(new_n5064));
  nor2 g04871(.a(new_n5064), .b(new_n4746), .O(new_n5065));
  inv1 g04872(.a(new_n5064), .O(new_n5066));
  nor2 g04873(.a(new_n5066), .b(new_n4745), .O(new_n5067));
  nor2 g04874(.a(new_n5067), .b(new_n5065), .O(new_n5068));
  nor2 g04875(.a(new_n5068), .b(new_n5057), .O(new_n5069));
  inv1 g04876(.a(new_n5057), .O(new_n5070));
  inv1 g04877(.a(new_n5068), .O(new_n5071));
  nor2 g04878(.a(new_n5071), .b(new_n5070), .O(new_n5072));
  nor2 g04879(.a(new_n5072), .b(new_n5069), .O(new_n5073));
  inv1 g04880(.a(new_n5073), .O(new_n5074));
  nor2 g04881(.a(new_n2826), .b(new_n438), .O(new_n5075));
  inv1 g04882(.a(new_n5075), .O(new_n5076));
  nor2 g04883(.a(new_n3533), .b(new_n295), .O(new_n5077));
  nor2 g04884(.a(new_n5077), .b(new_n4529), .O(new_n5078));
  inv1 g04885(.a(new_n4527), .O(new_n5079));
  nor2 g04886(.a(new_n3533), .b(new_n363), .O(new_n5080));
  inv1 g04887(.a(new_n5080), .O(new_n5081));
  nor2 g04888(.a(new_n5081), .b(new_n5079), .O(new_n5082));
  nor2 g04889(.a(new_n5082), .b(new_n5078), .O(new_n5083));
  nor2 g04890(.a(new_n5083), .b(new_n5076), .O(new_n5084));
  inv1 g04891(.a(new_n5083), .O(new_n5085));
  nor2 g04892(.a(new_n5085), .b(new_n5075), .O(new_n5086));
  nor2 g04893(.a(new_n5086), .b(new_n5084), .O(new_n5087));
  nor2 g04894(.a(new_n5087), .b(new_n5074), .O(new_n5088));
  inv1 g04895(.a(new_n5087), .O(new_n5089));
  nor2 g04896(.a(new_n5089), .b(new_n5073), .O(new_n5090));
  nor2 g04897(.a(new_n5090), .b(new_n5088), .O(new_n5091));
  nor2 g04898(.a(new_n5091), .b(new_n5044), .O(new_n5092));
  inv1 g04899(.a(new_n5044), .O(new_n5093));
  inv1 g04900(.a(new_n5091), .O(new_n5094));
  nor2 g04901(.a(new_n5094), .b(new_n5093), .O(new_n5095));
  nor2 g04902(.a(new_n5095), .b(new_n5092), .O(new_n5096));
  inv1 g04903(.a(new_n5096), .O(new_n5097));
  nor2 g04904(.a(new_n5097), .b(new_n5001), .O(new_n5098));
  inv1 g04905(.a(new_n5001), .O(new_n5099));
  nor2 g04906(.a(new_n5096), .b(new_n5099), .O(new_n5100));
  nor2 g04907(.a(new_n5100), .b(new_n5098), .O(new_n5101));
  inv1 g04908(.a(new_n5101), .O(new_n5102));
  nor2 g04909(.a(new_n5102), .b(new_n5000), .O(new_n5103));
  nor2 g04910(.a(new_n5101), .b(new_n4999), .O(new_n5104));
  nor2 g04911(.a(new_n5104), .b(new_n5103), .O(new_n5105));
  inv1 g04912(.a(new_n5105), .O(new_n5106));
  nor2 g04913(.a(new_n5106), .b(new_n4938), .O(new_n5107));
  nor2 g04914(.a(new_n5105), .b(new_n4937), .O(new_n5108));
  nor2 g04915(.a(new_n5108), .b(new_n5107), .O(new_n5109));
  nor2 g04916(.a(new_n5109), .b(new_n4879), .O(new_n5110));
  inv1 g04917(.a(new_n5109), .O(new_n5111));
  nor2 g04918(.a(new_n5111), .b(new_n4878), .O(new_n5112));
  nor2 g04919(.a(new_n5112), .b(new_n5110), .O(new_n5113));
  inv1 g04920(.a(new_n5113), .O(new_n5114));
  nor2 g04921(.a(new_n4873), .b(new_n4869), .O(new_n5115));
  nor2 g04922(.a(new_n5115), .b(new_n5114), .O(new_n5116));
  inv1 g04923(.a(new_n5115), .O(new_n5117));
  nor2 g04924(.a(new_n5117), .b(new_n5113), .O(new_n5118));
  nor2 g04925(.a(new_n5118), .b(new_n5116), .O(new_n5119));
  inv1 g04926(.a(new_n5119), .O(\asquared[42] ));
  nor2 g04927(.a(new_n5107), .b(new_n4936), .O(new_n5121));
  nor2 g04928(.a(new_n5103), .b(new_n5098), .O(new_n5122));
  nor2 g04929(.a(new_n4998), .b(new_n4991), .O(new_n5123));
  nor2 g04930(.a(new_n4894), .b(new_n4888), .O(new_n5124));
  inv1 g04931(.a(new_n5124), .O(new_n5125));
  nor2 g04932(.a(new_n4986), .b(new_n4969), .O(new_n5126));
  inv1 g04933(.a(new_n5126), .O(new_n5127));
  nor2 g04934(.a(new_n5127), .b(new_n5125), .O(new_n5128));
  nor2 g04935(.a(new_n5126), .b(new_n5124), .O(new_n5129));
  nor2 g04936(.a(new_n5129), .b(new_n5128), .O(new_n5130));
  nor2 g04937(.a(new_n5088), .b(new_n5069), .O(new_n5131));
  inv1 g04938(.a(new_n5131), .O(new_n5132));
  nor2 g04939(.a(new_n5132), .b(new_n5130), .O(new_n5133));
  inv1 g04940(.a(new_n5130), .O(new_n5134));
  nor2 g04941(.a(new_n5131), .b(new_n5134), .O(new_n5135));
  nor2 g04942(.a(new_n5135), .b(new_n5133), .O(new_n5136));
  inv1 g04943(.a(new_n5136), .O(new_n5137));
  nor2 g04944(.a(new_n5095), .b(new_n5043), .O(new_n5138));
  nor2 g04945(.a(new_n5138), .b(new_n5137), .O(new_n5139));
  inv1 g04946(.a(new_n5138), .O(new_n5140));
  nor2 g04947(.a(new_n5140), .b(new_n5136), .O(new_n5141));
  nor2 g04948(.a(new_n5141), .b(new_n5139), .O(new_n5142));
  inv1 g04949(.a(new_n5142), .O(new_n5143));
  nor2 g04950(.a(new_n5143), .b(new_n5123), .O(new_n5144));
  inv1 g04951(.a(new_n5123), .O(new_n5145));
  nor2 g04952(.a(new_n5142), .b(new_n5145), .O(new_n5146));
  nor2 g04953(.a(new_n5146), .b(new_n5144), .O(new_n5147));
  inv1 g04954(.a(new_n5147), .O(new_n5148));
  nor2 g04955(.a(new_n5148), .b(new_n5122), .O(new_n5149));
  inv1 g04956(.a(new_n5122), .O(new_n5150));
  nor2 g04957(.a(new_n5147), .b(new_n5150), .O(new_n5151));
  nor2 g04958(.a(new_n5151), .b(new_n5149), .O(new_n5152));
  inv1 g04959(.a(new_n5152), .O(new_n5153));
  nor2 g04960(.a(new_n4916), .b(new_n4911), .O(new_n5154));
  inv1 g04961(.a(new_n5154), .O(new_n5155));
  nor2 g04962(.a(new_n2506), .b(new_n613), .O(new_n5156));
  inv1 g04963(.a(new_n5156), .O(new_n5157));
  nor2 g04964(.a(new_n4093), .b(new_n229), .O(new_n5158));
  nor2 g04965(.a(new_n2660), .b(new_n569), .O(new_n5159));
  nor2 g04966(.a(new_n5159), .b(new_n5158), .O(new_n5160));
  inv1 g04967(.a(new_n5158), .O(new_n5161));
  inv1 g04968(.a(new_n5159), .O(new_n5162));
  nor2 g04969(.a(new_n5162), .b(new_n5161), .O(new_n5163));
  nor2 g04970(.a(new_n5163), .b(new_n5160), .O(new_n5164));
  nor2 g04971(.a(new_n5164), .b(new_n5157), .O(new_n5165));
  inv1 g04972(.a(new_n5164), .O(new_n5166));
  nor2 g04973(.a(new_n5166), .b(new_n5156), .O(new_n5167));
  nor2 g04974(.a(new_n5167), .b(new_n5165), .O(new_n5168));
  nor2 g04975(.a(new_n1493), .b(new_n1297), .O(new_n5169));
  nor2 g04976(.a(new_n4954), .b(new_n194), .O(new_n5170));
  nor2 g04977(.a(new_n5170), .b(new_n5169), .O(new_n5171));
  inv1 g04978(.a(new_n5169), .O(new_n5172));
  inv1 g04979(.a(new_n5170), .O(new_n5173));
  nor2 g04980(.a(new_n5173), .b(new_n5172), .O(new_n5174));
  nor2 g04981(.a(new_n5174), .b(new_n5171), .O(new_n5175));
  inv1 g04982(.a(new_n5175), .O(new_n5176));
  inv1 g04983(.a(new_n4903), .O(new_n5177));
  inv1 g04984(.a(\a[42] ), .O(new_n5178));
  nor2 g04985(.a(new_n5178), .b(new_n198), .O(new_n5179));
  inv1 g04986(.a(new_n5179), .O(new_n5180));
  nor2 g04987(.a(new_n5180), .b(new_n5177), .O(new_n5181));
  nor2 g04988(.a(new_n5179), .b(new_n4903), .O(new_n5182));
  nor2 g04989(.a(new_n5182), .b(new_n5181), .O(new_n5183));
  inv1 g04990(.a(new_n5183), .O(new_n5184));
  nor2 g04991(.a(new_n5184), .b(new_n5176), .O(new_n5185));
  nor2 g04992(.a(new_n5183), .b(new_n5175), .O(new_n5186));
  nor2 g04993(.a(new_n5186), .b(new_n5185), .O(new_n5187));
  inv1 g04994(.a(new_n5187), .O(new_n5188));
  nor2 g04995(.a(new_n5188), .b(new_n5168), .O(new_n5189));
  inv1 g04996(.a(new_n5168), .O(new_n5190));
  nor2 g04997(.a(new_n5187), .b(new_n5190), .O(new_n5191));
  nor2 g04998(.a(new_n5191), .b(new_n5189), .O(new_n5192));
  nor2 g04999(.a(new_n5192), .b(new_n5155), .O(new_n5193));
  inv1 g05000(.a(new_n5192), .O(new_n5194));
  nor2 g05001(.a(new_n5194), .b(new_n5154), .O(new_n5195));
  nor2 g05002(.a(new_n5195), .b(new_n5193), .O(new_n5196));
  nor2 g05003(.a(new_n4920), .b(new_n4900), .O(new_n5197));
  inv1 g05004(.a(new_n5197), .O(new_n5198));
  nor2 g05005(.a(new_n5198), .b(new_n5196), .O(new_n5199));
  inv1 g05006(.a(new_n5196), .O(new_n5200));
  nor2 g05007(.a(new_n5197), .b(new_n5200), .O(new_n5201));
  nor2 g05008(.a(new_n5201), .b(new_n5199), .O(new_n5202));
  inv1 g05009(.a(new_n5202), .O(new_n5203));
  nor2 g05010(.a(new_n5028), .b(new_n5021), .O(new_n5204));
  nor2 g05011(.a(new_n5067), .b(new_n5060), .O(new_n5205));
  nor2 g05012(.a(new_n5205), .b(new_n5204), .O(new_n5206));
  inv1 g05013(.a(new_n5204), .O(new_n5207));
  inv1 g05014(.a(new_n5205), .O(new_n5208));
  nor2 g05015(.a(new_n5208), .b(new_n5207), .O(new_n5209));
  nor2 g05016(.a(new_n5209), .b(new_n5206), .O(new_n5210));
  nor2 g05017(.a(new_n5013), .b(new_n5007), .O(new_n5211));
  nor2 g05018(.a(new_n5211), .b(new_n5210), .O(new_n5212));
  inv1 g05019(.a(new_n5210), .O(new_n5213));
  inv1 g05020(.a(new_n5211), .O(new_n5214));
  nor2 g05021(.a(new_n5214), .b(new_n5213), .O(new_n5215));
  nor2 g05022(.a(new_n5215), .b(new_n5212), .O(new_n5216));
  nor2 g05023(.a(new_n5037), .b(new_n5030), .O(new_n5217));
  inv1 g05024(.a(new_n5217), .O(new_n5218));
  nor2 g05025(.a(new_n5218), .b(new_n5216), .O(new_n5219));
  inv1 g05026(.a(new_n5216), .O(new_n5220));
  nor2 g05027(.a(new_n5217), .b(new_n5220), .O(new_n5221));
  nor2 g05028(.a(new_n5221), .b(new_n5219), .O(new_n5222));
  inv1 g05029(.a(new_n5222), .O(new_n5223));
  nor2 g05030(.a(new_n4984), .b(new_n4977), .O(new_n5224));
  nor2 g05031(.a(new_n5056), .b(new_n5048), .O(new_n5225));
  nor2 g05032(.a(new_n5225), .b(new_n5224), .O(new_n5226));
  inv1 g05033(.a(new_n5224), .O(new_n5227));
  inv1 g05034(.a(new_n5225), .O(new_n5228));
  nor2 g05035(.a(new_n5228), .b(new_n5227), .O(new_n5229));
  nor2 g05036(.a(new_n5229), .b(new_n5226), .O(new_n5230));
  nor2 g05037(.a(new_n4963), .b(new_n4960), .O(new_n5231));
  inv1 g05038(.a(new_n5231), .O(new_n5232));
  nor2 g05039(.a(new_n5232), .b(new_n5230), .O(new_n5233));
  inv1 g05040(.a(new_n5230), .O(new_n5234));
  nor2 g05041(.a(new_n5231), .b(new_n5234), .O(new_n5235));
  nor2 g05042(.a(new_n5235), .b(new_n5233), .O(new_n5236));
  inv1 g05043(.a(new_n5236), .O(new_n5237));
  nor2 g05044(.a(new_n5237), .b(new_n5223), .O(new_n5238));
  nor2 g05045(.a(new_n5236), .b(new_n5222), .O(new_n5239));
  nor2 g05046(.a(new_n5239), .b(new_n5238), .O(new_n5240));
  inv1 g05047(.a(new_n5240), .O(new_n5241));
  nor2 g05048(.a(new_n5241), .b(new_n5203), .O(new_n5242));
  nor2 g05049(.a(new_n5240), .b(new_n5202), .O(new_n5243));
  nor2 g05050(.a(new_n5243), .b(new_n5242), .O(new_n5244));
  inv1 g05051(.a(new_n5244), .O(new_n5245));
  nor2 g05052(.a(new_n4930), .b(new_n4924), .O(new_n5246));
  nor2 g05053(.a(new_n4950), .b(new_n4944), .O(new_n5247));
  inv1 g05054(.a(new_n5247), .O(new_n5248));
  nor2 g05055(.a(new_n3231), .b(new_n363), .O(new_n5249));
  nor2 g05056(.a(new_n3533), .b(new_n322), .O(new_n5250));
  nor2 g05057(.a(new_n5250), .b(new_n5249), .O(new_n5251));
  nor2 g05058(.a(new_n5081), .b(new_n5018), .O(new_n5252));
  nor2 g05059(.a(new_n5252), .b(new_n5251), .O(new_n5253));
  nor2 g05060(.a(new_n5253), .b(new_n4049), .O(new_n5254));
  inv1 g05061(.a(new_n5253), .O(new_n5255));
  nor2 g05062(.a(new_n5255), .b(new_n4048), .O(new_n5256));
  nor2 g05063(.a(new_n5256), .b(new_n5254), .O(new_n5257));
  nor2 g05064(.a(new_n3870), .b(new_n257), .O(new_n5258));
  inv1 g05065(.a(new_n5258), .O(new_n5259));
  nor2 g05066(.a(new_n3722), .b(new_n295), .O(new_n5260));
  nor2 g05067(.a(new_n2826), .b(new_n502), .O(new_n5261));
  nor2 g05068(.a(new_n5261), .b(new_n5260), .O(new_n5262));
  inv1 g05069(.a(new_n5260), .O(new_n5263));
  inv1 g05070(.a(new_n5261), .O(new_n5264));
  nor2 g05071(.a(new_n5264), .b(new_n5263), .O(new_n5265));
  nor2 g05072(.a(new_n5265), .b(new_n5262), .O(new_n5266));
  nor2 g05073(.a(new_n5266), .b(new_n5259), .O(new_n5267));
  inv1 g05074(.a(new_n5266), .O(new_n5268));
  nor2 g05075(.a(new_n5268), .b(new_n5258), .O(new_n5269));
  nor2 g05076(.a(new_n5269), .b(new_n5267), .O(new_n5270));
  nor2 g05077(.a(new_n5086), .b(new_n5078), .O(new_n5271));
  inv1 g05078(.a(new_n5271), .O(new_n5272));
  nor2 g05079(.a(new_n5272), .b(new_n5270), .O(new_n5273));
  inv1 g05080(.a(new_n5270), .O(new_n5274));
  nor2 g05081(.a(new_n5271), .b(new_n5274), .O(new_n5275));
  nor2 g05082(.a(new_n5275), .b(new_n5273), .O(new_n5276));
  inv1 g05083(.a(new_n5276), .O(new_n5277));
  nor2 g05084(.a(new_n5277), .b(new_n5257), .O(new_n5278));
  inv1 g05085(.a(new_n5257), .O(new_n5279));
  nor2 g05086(.a(new_n5276), .b(new_n5279), .O(new_n5280));
  nor2 g05087(.a(new_n5280), .b(new_n5278), .O(new_n5281));
  nor2 g05088(.a(new_n5281), .b(new_n5248), .O(new_n5282));
  inv1 g05089(.a(new_n5281), .O(new_n5283));
  nor2 g05090(.a(new_n5283), .b(new_n5247), .O(new_n5284));
  nor2 g05091(.a(new_n5284), .b(new_n5282), .O(new_n5285));
  inv1 g05092(.a(new_n5285), .O(new_n5286));
  nor2 g05093(.a(new_n2184), .b(new_n800), .O(new_n5287));
  inv1 g05094(.a(new_n5287), .O(new_n5288));
  nor2 g05095(.a(new_n4366), .b(new_n214), .O(new_n5289));
  nor2 g05096(.a(new_n2433), .b(new_n699), .O(new_n5290));
  nor2 g05097(.a(new_n5290), .b(new_n5289), .O(new_n5291));
  nor2 g05098(.a(new_n4366), .b(new_n699), .O(new_n5292));
  inv1 g05099(.a(new_n5292), .O(new_n5293));
  nor2 g05100(.a(new_n5293), .b(new_n2868), .O(new_n5294));
  nor2 g05101(.a(new_n5294), .b(new_n5291), .O(new_n5295));
  nor2 g05102(.a(new_n5295), .b(new_n5288), .O(new_n5296));
  inv1 g05103(.a(new_n5295), .O(new_n5297));
  nor2 g05104(.a(new_n5297), .b(new_n5287), .O(new_n5298));
  nor2 g05105(.a(new_n5298), .b(new_n5296), .O(new_n5299));
  inv1 g05106(.a(new_n5299), .O(new_n5300));
  nor2 g05107(.a(new_n1903), .b(new_n941), .O(new_n5301));
  inv1 g05108(.a(new_n5301), .O(new_n5302));
  nor2 g05109(.a(new_n1647), .b(new_n1199), .O(new_n5303));
  nor2 g05110(.a(new_n5303), .b(new_n5050), .O(new_n5304));
  inv1 g05111(.a(new_n5047), .O(new_n5305));
  nor2 g05112(.a(new_n1736), .b(new_n1199), .O(new_n5306));
  inv1 g05113(.a(new_n5306), .O(new_n5307));
  nor2 g05114(.a(new_n5307), .b(new_n5305), .O(new_n5308));
  nor2 g05115(.a(new_n5308), .b(new_n5304), .O(new_n5309));
  nor2 g05116(.a(new_n5309), .b(new_n5302), .O(new_n5310));
  inv1 g05117(.a(new_n5309), .O(new_n5311));
  nor2 g05118(.a(new_n5311), .b(new_n5301), .O(new_n5312));
  nor2 g05119(.a(new_n5312), .b(new_n5310), .O(new_n5313));
  nor2 g05120(.a(new_n4425), .b(new_n203), .O(new_n5314));
  nor2 g05121(.a(new_n2121), .b(new_n847), .O(new_n5315));
  nor2 g05122(.a(new_n5315), .b(new_n5314), .O(new_n5316));
  inv1 g05123(.a(new_n5314), .O(new_n5317));
  inv1 g05124(.a(new_n5315), .O(new_n5318));
  nor2 g05125(.a(new_n5318), .b(new_n5317), .O(new_n5319));
  nor2 g05126(.a(new_n5319), .b(new_n5316), .O(new_n5320));
  nor2 g05127(.a(new_n5320), .b(new_n4687), .O(new_n5321));
  inv1 g05128(.a(new_n5320), .O(new_n5322));
  nor2 g05129(.a(new_n5322), .b(new_n4686), .O(new_n5323));
  nor2 g05130(.a(new_n5323), .b(new_n5321), .O(new_n5324));
  nor2 g05131(.a(new_n5324), .b(new_n5313), .O(new_n5325));
  inv1 g05132(.a(new_n5313), .O(new_n5326));
  inv1 g05133(.a(new_n5324), .O(new_n5327));
  nor2 g05134(.a(new_n5327), .b(new_n5326), .O(new_n5328));
  nor2 g05135(.a(new_n5328), .b(new_n5325), .O(new_n5329));
  nor2 g05136(.a(new_n5329), .b(new_n5300), .O(new_n5330));
  inv1 g05137(.a(new_n5329), .O(new_n5331));
  nor2 g05138(.a(new_n5331), .b(new_n5299), .O(new_n5332));
  nor2 g05139(.a(new_n5332), .b(new_n5330), .O(new_n5333));
  inv1 g05140(.a(new_n5333), .O(new_n5334));
  nor2 g05141(.a(new_n5334), .b(new_n5286), .O(new_n5335));
  nor2 g05142(.a(new_n5333), .b(new_n5285), .O(new_n5336));
  nor2 g05143(.a(new_n5336), .b(new_n5335), .O(new_n5337));
  inv1 g05144(.a(new_n5337), .O(new_n5338));
  nor2 g05145(.a(new_n5338), .b(new_n5246), .O(new_n5339));
  inv1 g05146(.a(new_n5246), .O(new_n5340));
  nor2 g05147(.a(new_n5337), .b(new_n5340), .O(new_n5341));
  nor2 g05148(.a(new_n5341), .b(new_n5339), .O(new_n5342));
  inv1 g05149(.a(new_n5342), .O(new_n5343));
  nor2 g05150(.a(new_n5343), .b(new_n5245), .O(new_n5344));
  nor2 g05151(.a(new_n5342), .b(new_n5244), .O(new_n5345));
  nor2 g05152(.a(new_n5345), .b(new_n5344), .O(new_n5346));
  inv1 g05153(.a(new_n5346), .O(new_n5347));
  nor2 g05154(.a(new_n5347), .b(new_n5153), .O(new_n5348));
  nor2 g05155(.a(new_n5346), .b(new_n5152), .O(new_n5349));
  nor2 g05156(.a(new_n5349), .b(new_n5348), .O(new_n5350));
  inv1 g05157(.a(new_n5350), .O(new_n5351));
  nor2 g05158(.a(new_n5351), .b(new_n5121), .O(new_n5352));
  inv1 g05159(.a(new_n5121), .O(new_n5353));
  nor2 g05160(.a(new_n5350), .b(new_n5353), .O(new_n5354));
  nor2 g05161(.a(new_n5354), .b(new_n5352), .O(new_n5355));
  inv1 g05162(.a(new_n5355), .O(new_n5356));
  nor2 g05163(.a(new_n5116), .b(new_n5110), .O(new_n5357));
  nor2 g05164(.a(new_n5357), .b(new_n5356), .O(new_n5358));
  inv1 g05165(.a(new_n5357), .O(new_n5359));
  nor2 g05166(.a(new_n5359), .b(new_n5355), .O(new_n5360));
  nor2 g05167(.a(new_n5360), .b(new_n5358), .O(new_n5361));
  inv1 g05168(.a(new_n5361), .O(\asquared[43] ));
  nor2 g05169(.a(new_n5348), .b(new_n5149), .O(new_n5363));
  nor2 g05170(.a(new_n5144), .b(new_n5139), .O(new_n5364));
  nor2 g05171(.a(new_n5135), .b(new_n5129), .O(new_n5365));
  nor2 g05172(.a(new_n2121), .b(new_n941), .O(new_n5366));
  inv1 g05173(.a(new_n5366), .O(new_n5367));
  nor2 g05174(.a(new_n1903), .b(new_n1086), .O(new_n5368));
  nor2 g05175(.a(new_n5368), .b(new_n5306), .O(new_n5369));
  nor2 g05176(.a(new_n1903), .b(new_n1199), .O(new_n5370));
  inv1 g05177(.a(new_n5370), .O(new_n5371));
  nor2 g05178(.a(new_n5371), .b(new_n5051), .O(new_n5372));
  nor2 g05179(.a(new_n5372), .b(new_n5369), .O(new_n5373));
  nor2 g05180(.a(new_n5373), .b(new_n5367), .O(new_n5374));
  inv1 g05181(.a(new_n5373), .O(new_n5375));
  nor2 g05182(.a(new_n5375), .b(new_n5366), .O(new_n5376));
  nor2 g05183(.a(new_n5376), .b(new_n5374), .O(new_n5377));
  inv1 g05184(.a(new_n5377), .O(new_n5378));
  nor2 g05185(.a(new_n2506), .b(new_n699), .O(new_n5379));
  inv1 g05186(.a(new_n5379), .O(new_n5380));
  nor2 g05187(.a(new_n2184), .b(new_n847), .O(new_n5381));
  nor2 g05188(.a(new_n5381), .b(new_n4978), .O(new_n5382));
  nor2 g05189(.a(new_n2433), .b(new_n847), .O(new_n5383));
  inv1 g05190(.a(new_n5383), .O(new_n5384));
  nor2 g05191(.a(new_n5384), .b(new_n5288), .O(new_n5385));
  nor2 g05192(.a(new_n5385), .b(new_n5382), .O(new_n5386));
  nor2 g05193(.a(new_n5386), .b(new_n5380), .O(new_n5387));
  inv1 g05194(.a(new_n5386), .O(new_n5388));
  nor2 g05195(.a(new_n5388), .b(new_n5379), .O(new_n5389));
  nor2 g05196(.a(new_n5389), .b(new_n5387), .O(new_n5390));
  nor2 g05197(.a(new_n4425), .b(new_n214), .O(new_n5391));
  inv1 g05198(.a(new_n5391), .O(new_n5392));
  inv1 g05199(.a(\a[43] ), .O(new_n5393));
  nor2 g05200(.a(new_n5393), .b(new_n198), .O(new_n5394));
  nor2 g05201(.a(new_n4682), .b(new_n203), .O(new_n5395));
  nor2 g05202(.a(new_n5395), .b(new_n5394), .O(new_n5396));
  inv1 g05203(.a(new_n5394), .O(new_n5397));
  inv1 g05204(.a(new_n5395), .O(new_n5398));
  nor2 g05205(.a(new_n5398), .b(new_n5397), .O(new_n5399));
  nor2 g05206(.a(new_n5399), .b(new_n5396), .O(new_n5400));
  nor2 g05207(.a(new_n5400), .b(new_n5392), .O(new_n5401));
  inv1 g05208(.a(new_n5400), .O(new_n5402));
  nor2 g05209(.a(new_n5402), .b(new_n5391), .O(new_n5403));
  nor2 g05210(.a(new_n5403), .b(new_n5401), .O(new_n5404));
  nor2 g05211(.a(new_n5404), .b(new_n5390), .O(new_n5405));
  inv1 g05212(.a(new_n5390), .O(new_n5406));
  inv1 g05213(.a(new_n5404), .O(new_n5407));
  nor2 g05214(.a(new_n5407), .b(new_n5406), .O(new_n5408));
  nor2 g05215(.a(new_n5408), .b(new_n5405), .O(new_n5409));
  nor2 g05216(.a(new_n5409), .b(new_n5378), .O(new_n5410));
  inv1 g05217(.a(new_n5409), .O(new_n5411));
  nor2 g05218(.a(new_n5411), .b(new_n5377), .O(new_n5412));
  nor2 g05219(.a(new_n5412), .b(new_n5410), .O(new_n5413));
  inv1 g05220(.a(new_n5413), .O(new_n5414));
  nor2 g05221(.a(new_n4366), .b(new_n229), .O(new_n5415));
  nor2 g05222(.a(new_n2660), .b(new_n613), .O(new_n5416));
  nor2 g05223(.a(new_n5416), .b(new_n5415), .O(new_n5417));
  inv1 g05224(.a(new_n5415), .O(new_n5418));
  inv1 g05225(.a(new_n5416), .O(new_n5419));
  nor2 g05226(.a(new_n5419), .b(new_n5418), .O(new_n5420));
  nor2 g05227(.a(new_n5420), .b(new_n5417), .O(new_n5421));
  nor2 g05228(.a(new_n5421), .b(new_n4959), .O(new_n5422));
  inv1 g05229(.a(new_n5421), .O(new_n5423));
  nor2 g05230(.a(new_n5423), .b(new_n4958), .O(new_n5424));
  nor2 g05231(.a(new_n5424), .b(new_n5422), .O(new_n5425));
  inv1 g05232(.a(new_n5425), .O(new_n5426));
  nor2 g05233(.a(new_n3870), .b(new_n295), .O(new_n5427));
  nor2 g05234(.a(new_n3231), .b(new_n438), .O(new_n5428));
  nor2 g05235(.a(new_n3722), .b(new_n322), .O(new_n5429));
  nor2 g05236(.a(new_n5429), .b(new_n5428), .O(new_n5430));
  nor2 g05237(.a(new_n3722), .b(new_n438), .O(new_n5431));
  inv1 g05238(.a(new_n5431), .O(new_n5432));
  nor2 g05239(.a(new_n5432), .b(new_n5018), .O(new_n5433));
  nor2 g05240(.a(new_n5433), .b(new_n5430), .O(new_n5434));
  inv1 g05241(.a(new_n5434), .O(new_n5435));
  nor2 g05242(.a(new_n5435), .b(new_n5427), .O(new_n5436));
  inv1 g05243(.a(new_n5427), .O(new_n5437));
  nor2 g05244(.a(new_n5434), .b(new_n5437), .O(new_n5438));
  nor2 g05245(.a(new_n5438), .b(new_n5436), .O(new_n5439));
  nor2 g05246(.a(new_n1493), .b(new_n1425), .O(new_n5440));
  nor2 g05247(.a(new_n1647), .b(new_n1297), .O(new_n5441));
  nor2 g05248(.a(new_n5441), .b(new_n5440), .O(new_n5442));
  nor2 g05249(.a(new_n1647), .b(new_n1425), .O(new_n5443));
  inv1 g05250(.a(new_n5443), .O(new_n5444));
  nor2 g05251(.a(new_n5444), .b(new_n5172), .O(new_n5445));
  nor2 g05252(.a(new_n5445), .b(new_n5442), .O(new_n5446));
  nor2 g05253(.a(new_n5446), .b(new_n5081), .O(new_n5447));
  inv1 g05254(.a(new_n5446), .O(new_n5448));
  nor2 g05255(.a(new_n5448), .b(new_n5080), .O(new_n5449));
  nor2 g05256(.a(new_n5449), .b(new_n5447), .O(new_n5450));
  nor2 g05257(.a(new_n5450), .b(new_n5439), .O(new_n5451));
  inv1 g05258(.a(new_n5439), .O(new_n5452));
  inv1 g05259(.a(new_n5450), .O(new_n5453));
  nor2 g05260(.a(new_n5453), .b(new_n5452), .O(new_n5454));
  nor2 g05261(.a(new_n5454), .b(new_n5451), .O(new_n5455));
  nor2 g05262(.a(new_n5455), .b(new_n5426), .O(new_n5456));
  inv1 g05263(.a(new_n5455), .O(new_n5457));
  nor2 g05264(.a(new_n5457), .b(new_n5425), .O(new_n5458));
  nor2 g05265(.a(new_n5458), .b(new_n5456), .O(new_n5459));
  inv1 g05266(.a(new_n5459), .O(new_n5460));
  nor2 g05267(.a(new_n5460), .b(new_n5414), .O(new_n5461));
  nor2 g05268(.a(new_n5459), .b(new_n5413), .O(new_n5462));
  nor2 g05269(.a(new_n5462), .b(new_n5461), .O(new_n5463));
  inv1 g05270(.a(new_n5463), .O(new_n5464));
  nor2 g05271(.a(new_n5464), .b(new_n5365), .O(new_n5465));
  inv1 g05272(.a(new_n5365), .O(new_n5466));
  nor2 g05273(.a(new_n5463), .b(new_n5466), .O(new_n5467));
  nor2 g05274(.a(new_n5467), .b(new_n5465), .O(new_n5468));
  inv1 g05275(.a(new_n5468), .O(new_n5469));
  nor2 g05276(.a(new_n5469), .b(new_n5364), .O(new_n5470));
  inv1 g05277(.a(new_n5364), .O(new_n5471));
  nor2 g05278(.a(new_n5468), .b(new_n5471), .O(new_n5472));
  nor2 g05279(.a(new_n5472), .b(new_n5470), .O(new_n5473));
  inv1 g05280(.a(new_n5473), .O(new_n5474));
  nor2 g05281(.a(new_n5195), .b(new_n5189), .O(new_n5475));
  nor2 g05282(.a(new_n5269), .b(new_n5262), .O(new_n5476));
  nor2 g05283(.a(new_n5298), .b(new_n5291), .O(new_n5477));
  nor2 g05284(.a(new_n5477), .b(new_n5476), .O(new_n5478));
  inv1 g05285(.a(new_n5476), .O(new_n5479));
  inv1 g05286(.a(new_n5477), .O(new_n5480));
  nor2 g05287(.a(new_n5480), .b(new_n5479), .O(new_n5481));
  nor2 g05288(.a(new_n5481), .b(new_n5478), .O(new_n5482));
  nor2 g05289(.a(new_n5312), .b(new_n5304), .O(new_n5483));
  nor2 g05290(.a(new_n5483), .b(new_n5482), .O(new_n5484));
  inv1 g05291(.a(new_n5482), .O(new_n5485));
  inv1 g05292(.a(new_n5483), .O(new_n5486));
  nor2 g05293(.a(new_n5486), .b(new_n5485), .O(new_n5487));
  nor2 g05294(.a(new_n5487), .b(new_n5484), .O(new_n5488));
  nor2 g05295(.a(new_n5167), .b(new_n5160), .O(new_n5489));
  nor2 g05296(.a(new_n5323), .b(new_n5316), .O(new_n5490));
  nor2 g05297(.a(new_n5490), .b(new_n5489), .O(new_n5491));
  inv1 g05298(.a(new_n5489), .O(new_n5492));
  inv1 g05299(.a(new_n5490), .O(new_n5493));
  nor2 g05300(.a(new_n5493), .b(new_n5492), .O(new_n5494));
  nor2 g05301(.a(new_n5494), .b(new_n5491), .O(new_n5495));
  nor2 g05302(.a(new_n5185), .b(new_n5181), .O(new_n5496));
  inv1 g05303(.a(new_n5496), .O(new_n5497));
  nor2 g05304(.a(new_n5497), .b(new_n5495), .O(new_n5498));
  inv1 g05305(.a(new_n5495), .O(new_n5499));
  nor2 g05306(.a(new_n5496), .b(new_n5499), .O(new_n5500));
  nor2 g05307(.a(new_n5500), .b(new_n5498), .O(new_n5501));
  nor2 g05308(.a(new_n5501), .b(new_n5488), .O(new_n5502));
  inv1 g05309(.a(new_n5488), .O(new_n5503));
  inv1 g05310(.a(new_n5501), .O(new_n5504));
  nor2 g05311(.a(new_n5504), .b(new_n5503), .O(new_n5505));
  nor2 g05312(.a(new_n5505), .b(new_n5502), .O(new_n5506));
  inv1 g05313(.a(new_n5506), .O(new_n5507));
  nor2 g05314(.a(new_n5507), .b(new_n5475), .O(new_n5508));
  inv1 g05315(.a(new_n5475), .O(new_n5509));
  nor2 g05316(.a(new_n5506), .b(new_n5509), .O(new_n5510));
  nor2 g05317(.a(new_n5510), .b(new_n5508), .O(new_n5511));
  inv1 g05318(.a(new_n5511), .O(new_n5512));
  nor2 g05319(.a(new_n5235), .b(new_n5229), .O(new_n5513));
  inv1 g05320(.a(new_n5513), .O(new_n5514));
  nor2 g05321(.a(new_n5215), .b(new_n5209), .O(new_n5515));
  nor2 g05322(.a(new_n2826), .b(new_n569), .O(new_n5516));
  inv1 g05323(.a(new_n5516), .O(new_n5517));
  nor2 g05324(.a(new_n3057), .b(new_n502), .O(new_n5518));
  nor2 g05325(.a(new_n4093), .b(new_n257), .O(new_n5519));
  nor2 g05326(.a(new_n5519), .b(new_n5518), .O(new_n5520));
  inv1 g05327(.a(new_n5518), .O(new_n5521));
  inv1 g05328(.a(new_n5519), .O(new_n5522));
  nor2 g05329(.a(new_n5522), .b(new_n5521), .O(new_n5523));
  nor2 g05330(.a(new_n5523), .b(new_n5520), .O(new_n5524));
  nor2 g05331(.a(new_n5524), .b(new_n5517), .O(new_n5525));
  inv1 g05332(.a(new_n5524), .O(new_n5526));
  nor2 g05333(.a(new_n5526), .b(new_n5516), .O(new_n5527));
  nor2 g05334(.a(new_n5527), .b(new_n5525), .O(new_n5528));
  nor2 g05335(.a(new_n5528), .b(new_n5515), .O(new_n5529));
  inv1 g05336(.a(new_n5515), .O(new_n5530));
  inv1 g05337(.a(new_n5528), .O(new_n5531));
  nor2 g05338(.a(new_n5531), .b(new_n5530), .O(new_n5532));
  nor2 g05339(.a(new_n5532), .b(new_n5529), .O(new_n5533));
  nor2 g05340(.a(new_n5533), .b(new_n5514), .O(new_n5534));
  inv1 g05341(.a(new_n5533), .O(new_n5535));
  nor2 g05342(.a(new_n5535), .b(new_n5513), .O(new_n5536));
  nor2 g05343(.a(new_n5536), .b(new_n5534), .O(new_n5537));
  inv1 g05344(.a(new_n5537), .O(new_n5538));
  nor2 g05345(.a(new_n5238), .b(new_n5221), .O(new_n5539));
  nor2 g05346(.a(new_n5539), .b(new_n5538), .O(new_n5540));
  inv1 g05347(.a(new_n5539), .O(new_n5541));
  nor2 g05348(.a(new_n5541), .b(new_n5537), .O(new_n5542));
  nor2 g05349(.a(new_n5542), .b(new_n5540), .O(new_n5543));
  inv1 g05350(.a(new_n5543), .O(new_n5544));
  nor2 g05351(.a(new_n5544), .b(new_n5512), .O(new_n5545));
  nor2 g05352(.a(new_n5543), .b(new_n5511), .O(new_n5546));
  nor2 g05353(.a(new_n5546), .b(new_n5545), .O(new_n5547));
  inv1 g05354(.a(new_n5547), .O(new_n5548));
  nor2 g05355(.a(new_n5548), .b(new_n5474), .O(new_n5549));
  nor2 g05356(.a(new_n5547), .b(new_n5473), .O(new_n5550));
  nor2 g05357(.a(new_n5550), .b(new_n5549), .O(new_n5551));
  inv1 g05358(.a(new_n5551), .O(new_n5552));
  nor2 g05359(.a(new_n5344), .b(new_n5339), .O(new_n5553));
  nor2 g05360(.a(new_n5242), .b(new_n5201), .O(new_n5554));
  nor2 g05361(.a(new_n5335), .b(new_n5284), .O(new_n5555));
  nor2 g05362(.a(new_n5278), .b(new_n5273), .O(new_n5556));
  nor2 g05363(.a(new_n1692), .b(new_n5178), .O(new_n5557));
  nor2 g05364(.a(new_n5178), .b(new_n194), .O(new_n5558));
  nor2 g05365(.a(new_n5558), .b(\a[22] ), .O(new_n5559));
  nor2 g05366(.a(new_n5559), .b(new_n5557), .O(new_n5560));
  nor2 g05367(.a(new_n5560), .b(new_n5174), .O(new_n5561));
  inv1 g05368(.a(new_n5174), .O(new_n5562));
  nor2 g05369(.a(new_n5562), .b(\a[42] ), .O(new_n5563));
  nor2 g05370(.a(new_n5563), .b(new_n5561), .O(new_n5564));
  inv1 g05371(.a(new_n5564), .O(new_n5565));
  nor2 g05372(.a(new_n5256), .b(new_n5251), .O(new_n5566));
  inv1 g05373(.a(new_n5566), .O(new_n5567));
  nor2 g05374(.a(new_n5567), .b(new_n5565), .O(new_n5568));
  nor2 g05375(.a(new_n5566), .b(new_n5564), .O(new_n5569));
  nor2 g05376(.a(new_n5569), .b(new_n5568), .O(new_n5570));
  inv1 g05377(.a(new_n5570), .O(new_n5571));
  nor2 g05378(.a(new_n5571), .b(new_n5556), .O(new_n5572));
  inv1 g05379(.a(new_n5556), .O(new_n5573));
  nor2 g05380(.a(new_n5570), .b(new_n5573), .O(new_n5574));
  nor2 g05381(.a(new_n5574), .b(new_n5572), .O(new_n5575));
  inv1 g05382(.a(new_n5575), .O(new_n5576));
  nor2 g05383(.a(new_n5332), .b(new_n5325), .O(new_n5577));
  nor2 g05384(.a(new_n5577), .b(new_n5576), .O(new_n5578));
  inv1 g05385(.a(new_n5577), .O(new_n5579));
  nor2 g05386(.a(new_n5579), .b(new_n5575), .O(new_n5580));
  nor2 g05387(.a(new_n5580), .b(new_n5578), .O(new_n5581));
  inv1 g05388(.a(new_n5581), .O(new_n5582));
  nor2 g05389(.a(new_n5582), .b(new_n5555), .O(new_n5583));
  inv1 g05390(.a(new_n5555), .O(new_n5584));
  nor2 g05391(.a(new_n5581), .b(new_n5584), .O(new_n5585));
  nor2 g05392(.a(new_n5585), .b(new_n5583), .O(new_n5586));
  inv1 g05393(.a(new_n5586), .O(new_n5587));
  nor2 g05394(.a(new_n5587), .b(new_n5554), .O(new_n5588));
  inv1 g05395(.a(new_n5554), .O(new_n5589));
  nor2 g05396(.a(new_n5586), .b(new_n5589), .O(new_n5590));
  nor2 g05397(.a(new_n5590), .b(new_n5588), .O(new_n5591));
  inv1 g05398(.a(new_n5591), .O(new_n5592));
  nor2 g05399(.a(new_n5592), .b(new_n5553), .O(new_n5593));
  inv1 g05400(.a(new_n5553), .O(new_n5594));
  nor2 g05401(.a(new_n5591), .b(new_n5594), .O(new_n5595));
  nor2 g05402(.a(new_n5595), .b(new_n5593), .O(new_n5596));
  inv1 g05403(.a(new_n5596), .O(new_n5597));
  nor2 g05404(.a(new_n5597), .b(new_n5552), .O(new_n5598));
  nor2 g05405(.a(new_n5596), .b(new_n5551), .O(new_n5599));
  nor2 g05406(.a(new_n5599), .b(new_n5598), .O(new_n5600));
  inv1 g05407(.a(new_n5600), .O(new_n5601));
  nor2 g05408(.a(new_n5601), .b(new_n5363), .O(new_n5602));
  inv1 g05409(.a(new_n5363), .O(new_n5603));
  nor2 g05410(.a(new_n5600), .b(new_n5603), .O(new_n5604));
  nor2 g05411(.a(new_n5604), .b(new_n5602), .O(new_n5605));
  inv1 g05412(.a(new_n5605), .O(new_n5606));
  nor2 g05413(.a(new_n5358), .b(new_n5354), .O(new_n5607));
  nor2 g05414(.a(new_n5607), .b(new_n5606), .O(new_n5608));
  inv1 g05415(.a(new_n5607), .O(new_n5609));
  nor2 g05416(.a(new_n5609), .b(new_n5605), .O(new_n5610));
  nor2 g05417(.a(new_n5610), .b(new_n5608), .O(new_n5611));
  inv1 g05418(.a(new_n5611), .O(\asquared[44] ));
  nor2 g05419(.a(new_n5598), .b(new_n5593), .O(new_n5613));
  nor2 g05420(.a(new_n5549), .b(new_n5470), .O(new_n5614));
  nor2 g05421(.a(new_n5545), .b(new_n5540), .O(new_n5615));
  nor2 g05422(.a(new_n5465), .b(new_n5461), .O(new_n5616));
  nor2 g05423(.a(new_n5403), .b(new_n5396), .O(new_n5617));
  nor2 g05424(.a(new_n5424), .b(new_n5417), .O(new_n5618));
  nor2 g05425(.a(new_n5618), .b(new_n5617), .O(new_n5619));
  inv1 g05426(.a(new_n5617), .O(new_n5620));
  inv1 g05427(.a(new_n5618), .O(new_n5621));
  nor2 g05428(.a(new_n5621), .b(new_n5620), .O(new_n5622));
  nor2 g05429(.a(new_n5622), .b(new_n5619), .O(new_n5623));
  nor2 g05430(.a(new_n5376), .b(new_n5369), .O(new_n5624));
  nor2 g05431(.a(new_n5624), .b(new_n5623), .O(new_n5625));
  inv1 g05432(.a(new_n5623), .O(new_n5626));
  inv1 g05433(.a(new_n5624), .O(new_n5627));
  nor2 g05434(.a(new_n5627), .b(new_n5626), .O(new_n5628));
  nor2 g05435(.a(new_n5628), .b(new_n5625), .O(new_n5629));
  inv1 g05436(.a(new_n5629), .O(new_n5630));
  nor2 g05437(.a(new_n5412), .b(new_n5405), .O(new_n5631));
  inv1 g05438(.a(new_n5631), .O(new_n5632));
  nor2 g05439(.a(new_n5458), .b(new_n5451), .O(new_n5633));
  inv1 g05440(.a(new_n5633), .O(new_n5634));
  nor2 g05441(.a(new_n5634), .b(new_n5632), .O(new_n5635));
  nor2 g05442(.a(new_n5633), .b(new_n5631), .O(new_n5636));
  nor2 g05443(.a(new_n5636), .b(new_n5635), .O(new_n5637));
  inv1 g05444(.a(new_n5637), .O(new_n5638));
  nor2 g05445(.a(new_n5638), .b(new_n5630), .O(new_n5639));
  nor2 g05446(.a(new_n5637), .b(new_n5629), .O(new_n5640));
  nor2 g05447(.a(new_n5640), .b(new_n5639), .O(new_n5641));
  inv1 g05448(.a(new_n5641), .O(new_n5642));
  nor2 g05449(.a(new_n5642), .b(new_n5616), .O(new_n5643));
  inv1 g05450(.a(new_n5616), .O(new_n5644));
  nor2 g05451(.a(new_n5641), .b(new_n5644), .O(new_n5645));
  nor2 g05452(.a(new_n5645), .b(new_n5643), .O(new_n5646));
  inv1 g05453(.a(new_n5646), .O(new_n5647));
  nor2 g05454(.a(new_n5647), .b(new_n5615), .O(new_n5648));
  inv1 g05455(.a(new_n5615), .O(new_n5649));
  nor2 g05456(.a(new_n5646), .b(new_n5649), .O(new_n5650));
  nor2 g05457(.a(new_n5650), .b(new_n5648), .O(new_n5651));
  inv1 g05458(.a(new_n5651), .O(new_n5652));
  nor2 g05459(.a(new_n5652), .b(new_n5614), .O(new_n5653));
  inv1 g05460(.a(new_n5614), .O(new_n5654));
  nor2 g05461(.a(new_n5651), .b(new_n5654), .O(new_n5655));
  nor2 g05462(.a(new_n5655), .b(new_n5653), .O(new_n5656));
  inv1 g05463(.a(new_n5656), .O(new_n5657));
  nor2 g05464(.a(new_n5588), .b(new_n5583), .O(new_n5658));
  inv1 g05465(.a(new_n5658), .O(new_n5659));
  nor2 g05466(.a(new_n5578), .b(new_n5572), .O(new_n5660));
  nor2 g05467(.a(new_n4366), .b(new_n257), .O(new_n5661));
  inv1 g05468(.a(new_n5661), .O(new_n5662));
  nor2 g05469(.a(new_n4093), .b(new_n295), .O(new_n5663));
  nor2 g05470(.a(new_n5663), .b(new_n3235), .O(new_n5664));
  nor2 g05471(.a(new_n4093), .b(new_n502), .O(new_n5665));
  inv1 g05472(.a(new_n5665), .O(new_n5666));
  nor2 g05473(.a(new_n5666), .b(new_n4696), .O(new_n5667));
  nor2 g05474(.a(new_n5667), .b(new_n5664), .O(new_n5668));
  nor2 g05475(.a(new_n5668), .b(new_n5662), .O(new_n5669));
  inv1 g05476(.a(new_n5668), .O(new_n5670));
  nor2 g05477(.a(new_n5670), .b(new_n5661), .O(new_n5671));
  nor2 g05478(.a(new_n5671), .b(new_n5669), .O(new_n5672));
  inv1 g05479(.a(new_n5672), .O(new_n5673));
  nor2 g05480(.a(new_n4954), .b(new_n203), .O(new_n5674));
  nor2 g05481(.a(new_n2506), .b(new_n800), .O(new_n5675));
  nor2 g05482(.a(new_n2184), .b(new_n941), .O(new_n5676));
  nor2 g05483(.a(new_n5676), .b(new_n5675), .O(new_n5677));
  nor2 g05484(.a(new_n2506), .b(new_n941), .O(new_n5678));
  inv1 g05485(.a(new_n5678), .O(new_n5679));
  nor2 g05486(.a(new_n5679), .b(new_n5288), .O(new_n5680));
  nor2 g05487(.a(new_n5680), .b(new_n5677), .O(new_n5681));
  inv1 g05488(.a(new_n5681), .O(new_n5682));
  nor2 g05489(.a(new_n5682), .b(new_n5674), .O(new_n5683));
  inv1 g05490(.a(new_n5674), .O(new_n5684));
  nor2 g05491(.a(new_n5681), .b(new_n5684), .O(new_n5685));
  nor2 g05492(.a(new_n5685), .b(new_n5683), .O(new_n5686));
  nor2 g05493(.a(new_n2121), .b(new_n1086), .O(new_n5687));
  inv1 g05494(.a(new_n5687), .O(new_n5688));
  nor2 g05495(.a(new_n1736), .b(new_n1297), .O(new_n5689));
  nor2 g05496(.a(new_n5689), .b(new_n5370), .O(new_n5690));
  nor2 g05497(.a(new_n1903), .b(new_n1297), .O(new_n5691));
  inv1 g05498(.a(new_n5691), .O(new_n5692));
  nor2 g05499(.a(new_n5692), .b(new_n5307), .O(new_n5693));
  nor2 g05500(.a(new_n5693), .b(new_n5690), .O(new_n5694));
  nor2 g05501(.a(new_n5694), .b(new_n5688), .O(new_n5695));
  inv1 g05502(.a(new_n5694), .O(new_n5696));
  nor2 g05503(.a(new_n5696), .b(new_n5687), .O(new_n5697));
  nor2 g05504(.a(new_n5697), .b(new_n5695), .O(new_n5698));
  nor2 g05505(.a(new_n5698), .b(new_n5686), .O(new_n5699));
  inv1 g05506(.a(new_n5686), .O(new_n5700));
  inv1 g05507(.a(new_n5698), .O(new_n5701));
  nor2 g05508(.a(new_n5701), .b(new_n5700), .O(new_n5702));
  nor2 g05509(.a(new_n5702), .b(new_n5699), .O(new_n5703));
  nor2 g05510(.a(new_n5703), .b(new_n5673), .O(new_n5704));
  inv1 g05511(.a(new_n5703), .O(new_n5705));
  nor2 g05512(.a(new_n5705), .b(new_n5672), .O(new_n5706));
  nor2 g05513(.a(new_n5706), .b(new_n5704), .O(new_n5707));
  nor2 g05514(.a(new_n4425), .b(new_n229), .O(new_n5708));
  inv1 g05515(.a(new_n5708), .O(new_n5709));
  nor2 g05516(.a(new_n3057), .b(new_n569), .O(new_n5710));
  nor2 g05517(.a(new_n2826), .b(new_n613), .O(new_n5711));
  nor2 g05518(.a(new_n5711), .b(new_n5710), .O(new_n5712));
  nor2 g05519(.a(new_n3057), .b(new_n613), .O(new_n5713));
  inv1 g05520(.a(new_n5713), .O(new_n5714));
  nor2 g05521(.a(new_n5714), .b(new_n5517), .O(new_n5715));
  nor2 g05522(.a(new_n5715), .b(new_n5712), .O(new_n5716));
  nor2 g05523(.a(new_n5716), .b(new_n5709), .O(new_n5717));
  inv1 g05524(.a(new_n5716), .O(new_n5718));
  nor2 g05525(.a(new_n5718), .b(new_n5708), .O(new_n5719));
  nor2 g05526(.a(new_n5719), .b(new_n5717), .O(new_n5720));
  inv1 g05527(.a(new_n5720), .O(new_n5721));
  nor2 g05528(.a(new_n3870), .b(new_n322), .O(new_n5722));
  inv1 g05529(.a(new_n5722), .O(new_n5723));
  nor2 g05530(.a(new_n3722), .b(new_n363), .O(new_n5724));
  nor2 g05531(.a(new_n5724), .b(new_n4606), .O(new_n5725));
  nor2 g05532(.a(new_n5432), .b(new_n5081), .O(new_n5726));
  nor2 g05533(.a(new_n5726), .b(new_n5725), .O(new_n5727));
  nor2 g05534(.a(new_n5727), .b(new_n5723), .O(new_n5728));
  inv1 g05535(.a(new_n5727), .O(new_n5729));
  nor2 g05536(.a(new_n5729), .b(new_n5722), .O(new_n5730));
  nor2 g05537(.a(new_n5730), .b(new_n5728), .O(new_n5731));
  nor2 g05538(.a(new_n4682), .b(new_n214), .O(new_n5732));
  nor2 g05539(.a(new_n2660), .b(new_n699), .O(new_n5733));
  nor2 g05540(.a(new_n5733), .b(new_n5732), .O(new_n5734));
  inv1 g05541(.a(new_n5732), .O(new_n5735));
  inv1 g05542(.a(new_n5733), .O(new_n5736));
  nor2 g05543(.a(new_n5736), .b(new_n5735), .O(new_n5737));
  nor2 g05544(.a(new_n5737), .b(new_n5734), .O(new_n5738));
  nor2 g05545(.a(new_n5738), .b(new_n5384), .O(new_n5739));
  inv1 g05546(.a(new_n5738), .O(new_n5740));
  nor2 g05547(.a(new_n5740), .b(new_n5383), .O(new_n5741));
  nor2 g05548(.a(new_n5741), .b(new_n5739), .O(new_n5742));
  nor2 g05549(.a(new_n5742), .b(new_n5731), .O(new_n5743));
  inv1 g05550(.a(new_n5731), .O(new_n5744));
  inv1 g05551(.a(new_n5742), .O(new_n5745));
  nor2 g05552(.a(new_n5745), .b(new_n5744), .O(new_n5746));
  nor2 g05553(.a(new_n5746), .b(new_n5743), .O(new_n5747));
  nor2 g05554(.a(new_n5747), .b(new_n5721), .O(new_n5748));
  inv1 g05555(.a(new_n5747), .O(new_n5749));
  nor2 g05556(.a(new_n5749), .b(new_n5720), .O(new_n5750));
  nor2 g05557(.a(new_n5750), .b(new_n5748), .O(new_n5751));
  nor2 g05558(.a(new_n5751), .b(new_n5707), .O(new_n5752));
  inv1 g05559(.a(new_n5707), .O(new_n5753));
  inv1 g05560(.a(new_n5751), .O(new_n5754));
  nor2 g05561(.a(new_n5754), .b(new_n5753), .O(new_n5755));
  nor2 g05562(.a(new_n5755), .b(new_n5752), .O(new_n5756));
  inv1 g05563(.a(new_n5756), .O(new_n5757));
  nor2 g05564(.a(new_n5757), .b(new_n5660), .O(new_n5758));
  inv1 g05565(.a(new_n5660), .O(new_n5759));
  nor2 g05566(.a(new_n5756), .b(new_n5759), .O(new_n5760));
  nor2 g05567(.a(new_n5760), .b(new_n5758), .O(new_n5761));
  nor2 g05568(.a(new_n5761), .b(new_n5659), .O(new_n5762));
  inv1 g05569(.a(new_n5761), .O(new_n5763));
  nor2 g05570(.a(new_n5763), .b(new_n5658), .O(new_n5764));
  nor2 g05571(.a(new_n5764), .b(new_n5762), .O(new_n5765));
  inv1 g05572(.a(new_n5765), .O(new_n5766));
  nor2 g05573(.a(new_n5536), .b(new_n5529), .O(new_n5767));
  inv1 g05574(.a(new_n5767), .O(new_n5768));
  nor2 g05575(.a(new_n5393), .b(new_n194), .O(new_n5769));
  nor2 g05576(.a(new_n5769), .b(new_n5443), .O(new_n5770));
  inv1 g05577(.a(new_n5769), .O(new_n5771));
  nor2 g05578(.a(new_n5771), .b(new_n5444), .O(new_n5772));
  nor2 g05579(.a(new_n5772), .b(new_n5770), .O(new_n5773));
  nor2 g05580(.a(new_n5449), .b(new_n5442), .O(new_n5774));
  nor2 g05581(.a(new_n5774), .b(new_n5773), .O(new_n5775));
  inv1 g05582(.a(new_n5773), .O(new_n5776));
  inv1 g05583(.a(new_n5774), .O(new_n5777));
  nor2 g05584(.a(new_n5777), .b(new_n5776), .O(new_n5778));
  nor2 g05585(.a(new_n5778), .b(new_n5775), .O(new_n5779));
  inv1 g05586(.a(new_n5779), .O(new_n5780));
  nor2 g05587(.a(new_n5436), .b(new_n5430), .O(new_n5781));
  inv1 g05588(.a(new_n5781), .O(new_n5782));
  nor2 g05589(.a(new_n5782), .b(new_n5780), .O(new_n5783));
  nor2 g05590(.a(new_n5781), .b(new_n5779), .O(new_n5784));
  nor2 g05591(.a(new_n5784), .b(new_n5783), .O(new_n5785));
  inv1 g05592(.a(new_n5785), .O(new_n5786));
  nor2 g05593(.a(new_n5527), .b(new_n5520), .O(new_n5787));
  nor2 g05594(.a(new_n5389), .b(new_n5382), .O(new_n5788));
  nor2 g05595(.a(new_n5788), .b(new_n5787), .O(new_n5789));
  inv1 g05596(.a(new_n5787), .O(new_n5790));
  inv1 g05597(.a(new_n5788), .O(new_n5791));
  nor2 g05598(.a(new_n5791), .b(new_n5790), .O(new_n5792));
  nor2 g05599(.a(new_n5792), .b(new_n5789), .O(new_n5793));
  inv1 g05600(.a(new_n5793), .O(new_n5794));
  inv1 g05601(.a(new_n5557), .O(new_n5795));
  inv1 g05602(.a(\a[44] ), .O(new_n5796));
  nor2 g05603(.a(new_n5796), .b(new_n198), .O(new_n5797));
  nor2 g05604(.a(new_n5178), .b(new_n196), .O(new_n5798));
  nor2 g05605(.a(new_n5798), .b(new_n5797), .O(new_n5799));
  nor2 g05606(.a(new_n5796), .b(new_n196), .O(new_n5800));
  inv1 g05607(.a(new_n5800), .O(new_n5801));
  nor2 g05608(.a(new_n5801), .b(new_n5180), .O(new_n5802));
  nor2 g05609(.a(new_n5802), .b(new_n5799), .O(new_n5803));
  nor2 g05610(.a(new_n5803), .b(new_n5795), .O(new_n5804));
  inv1 g05611(.a(new_n5803), .O(new_n5805));
  nor2 g05612(.a(new_n5805), .b(new_n5557), .O(new_n5806));
  nor2 g05613(.a(new_n5806), .b(new_n5804), .O(new_n5807));
  nor2 g05614(.a(new_n5807), .b(new_n5794), .O(new_n5808));
  inv1 g05615(.a(new_n5807), .O(new_n5809));
  nor2 g05616(.a(new_n5809), .b(new_n5793), .O(new_n5810));
  nor2 g05617(.a(new_n5810), .b(new_n5808), .O(new_n5811));
  inv1 g05618(.a(new_n5811), .O(new_n5812));
  nor2 g05619(.a(new_n5812), .b(new_n5786), .O(new_n5813));
  nor2 g05620(.a(new_n5811), .b(new_n5785), .O(new_n5814));
  nor2 g05621(.a(new_n5814), .b(new_n5813), .O(new_n5815));
  nor2 g05622(.a(new_n5815), .b(new_n5768), .O(new_n5816));
  inv1 g05623(.a(new_n5815), .O(new_n5817));
  nor2 g05624(.a(new_n5817), .b(new_n5767), .O(new_n5818));
  nor2 g05625(.a(new_n5818), .b(new_n5816), .O(new_n5819));
  nor2 g05626(.a(new_n5508), .b(new_n5505), .O(new_n5820));
  nor2 g05627(.a(new_n5500), .b(new_n5494), .O(new_n5821));
  inv1 g05628(.a(new_n5821), .O(new_n5822));
  nor2 g05629(.a(new_n5568), .b(new_n5563), .O(new_n5823));
  inv1 g05630(.a(new_n5823), .O(new_n5824));
  nor2 g05631(.a(new_n5824), .b(new_n5822), .O(new_n5825));
  nor2 g05632(.a(new_n5823), .b(new_n5821), .O(new_n5826));
  nor2 g05633(.a(new_n5826), .b(new_n5825), .O(new_n5827));
  nor2 g05634(.a(new_n5487), .b(new_n5481), .O(new_n5828));
  inv1 g05635(.a(new_n5828), .O(new_n5829));
  nor2 g05636(.a(new_n5829), .b(new_n5827), .O(new_n5830));
  inv1 g05637(.a(new_n5827), .O(new_n5831));
  nor2 g05638(.a(new_n5828), .b(new_n5831), .O(new_n5832));
  nor2 g05639(.a(new_n5832), .b(new_n5830), .O(new_n5833));
  inv1 g05640(.a(new_n5833), .O(new_n5834));
  nor2 g05641(.a(new_n5834), .b(new_n5820), .O(new_n5835));
  inv1 g05642(.a(new_n5820), .O(new_n5836));
  nor2 g05643(.a(new_n5833), .b(new_n5836), .O(new_n5837));
  nor2 g05644(.a(new_n5837), .b(new_n5835), .O(new_n5838));
  nor2 g05645(.a(new_n5838), .b(new_n5819), .O(new_n5839));
  inv1 g05646(.a(new_n5819), .O(new_n5840));
  inv1 g05647(.a(new_n5838), .O(new_n5841));
  nor2 g05648(.a(new_n5841), .b(new_n5840), .O(new_n5842));
  nor2 g05649(.a(new_n5842), .b(new_n5839), .O(new_n5843));
  inv1 g05650(.a(new_n5843), .O(new_n5844));
  nor2 g05651(.a(new_n5844), .b(new_n5766), .O(new_n5845));
  nor2 g05652(.a(new_n5843), .b(new_n5765), .O(new_n5846));
  nor2 g05653(.a(new_n5846), .b(new_n5845), .O(new_n5847));
  inv1 g05654(.a(new_n5847), .O(new_n5848));
  nor2 g05655(.a(new_n5848), .b(new_n5657), .O(new_n5849));
  nor2 g05656(.a(new_n5847), .b(new_n5656), .O(new_n5850));
  nor2 g05657(.a(new_n5850), .b(new_n5849), .O(new_n5851));
  inv1 g05658(.a(new_n5851), .O(new_n5852));
  nor2 g05659(.a(new_n5852), .b(new_n5613), .O(new_n5853));
  inv1 g05660(.a(new_n5613), .O(new_n5854));
  nor2 g05661(.a(new_n5851), .b(new_n5854), .O(new_n5855));
  nor2 g05662(.a(new_n5855), .b(new_n5853), .O(new_n5856));
  inv1 g05663(.a(new_n5856), .O(new_n5857));
  nor2 g05664(.a(new_n5608), .b(new_n5604), .O(new_n5858));
  nor2 g05665(.a(new_n5858), .b(new_n5857), .O(new_n5859));
  inv1 g05666(.a(new_n5858), .O(new_n5860));
  nor2 g05667(.a(new_n5860), .b(new_n5856), .O(new_n5861));
  nor2 g05668(.a(new_n5861), .b(new_n5859), .O(new_n5862));
  inv1 g05669(.a(new_n5862), .O(\asquared[45] ));
  nor2 g05670(.a(new_n5849), .b(new_n5653), .O(new_n5864));
  nor2 g05671(.a(new_n5845), .b(new_n5764), .O(new_n5865));
  inv1 g05672(.a(new_n5865), .O(new_n5866));
  nor2 g05673(.a(new_n5806), .b(new_n5799), .O(new_n5867));
  nor2 g05674(.a(new_n5683), .b(new_n5677), .O(new_n5868));
  nor2 g05675(.a(new_n5868), .b(new_n5867), .O(new_n5869));
  inv1 g05676(.a(new_n5867), .O(new_n5870));
  inv1 g05677(.a(new_n5868), .O(new_n5871));
  nor2 g05678(.a(new_n5871), .b(new_n5870), .O(new_n5872));
  nor2 g05679(.a(new_n5872), .b(new_n5869), .O(new_n5873));
  nor2 g05680(.a(new_n5697), .b(new_n5690), .O(new_n5874));
  nor2 g05681(.a(new_n5874), .b(new_n5873), .O(new_n5875));
  inv1 g05682(.a(new_n5873), .O(new_n5876));
  inv1 g05683(.a(new_n5874), .O(new_n5877));
  nor2 g05684(.a(new_n5877), .b(new_n5876), .O(new_n5878));
  nor2 g05685(.a(new_n5878), .b(new_n5875), .O(new_n5879));
  nor2 g05686(.a(new_n5832), .b(new_n5826), .O(new_n5880));
  inv1 g05687(.a(new_n5880), .O(new_n5881));
  nor2 g05688(.a(new_n5881), .b(new_n5879), .O(new_n5882));
  inv1 g05689(.a(new_n5879), .O(new_n5883));
  nor2 g05690(.a(new_n5880), .b(new_n5883), .O(new_n5884));
  nor2 g05691(.a(new_n5884), .b(new_n5882), .O(new_n5885));
  inv1 g05692(.a(new_n5885), .O(new_n5886));
  nor2 g05693(.a(new_n5178), .b(new_n203), .O(new_n5887));
  nor2 g05694(.a(new_n5887), .b(new_n5772), .O(new_n5888));
  inv1 g05695(.a(new_n5772), .O(new_n5889));
  inv1 g05696(.a(new_n5887), .O(new_n5890));
  nor2 g05697(.a(new_n5890), .b(new_n5889), .O(new_n5891));
  nor2 g05698(.a(new_n5891), .b(new_n5888), .O(new_n5892));
  inv1 g05699(.a(new_n5892), .O(new_n5893));
  nor2 g05700(.a(new_n1745), .b(new_n5796), .O(new_n5894));
  nor2 g05701(.a(new_n5894), .b(new_n1647), .O(new_n5895));
  nor2 g05702(.a(\a[23] ), .b(new_n194), .O(new_n5896));
  inv1 g05703(.a(new_n5896), .O(new_n5897));
  nor2 g05704(.a(new_n5897), .b(new_n5796), .O(new_n5898));
  nor2 g05705(.a(new_n5898), .b(new_n5895), .O(new_n5899));
  nor2 g05706(.a(new_n5899), .b(new_n5893), .O(new_n5900));
  inv1 g05707(.a(new_n5899), .O(new_n5901));
  nor2 g05708(.a(new_n5901), .b(new_n5892), .O(new_n5902));
  nor2 g05709(.a(new_n5902), .b(new_n5900), .O(new_n5903));
  inv1 g05710(.a(new_n5903), .O(new_n5904));
  nor2 g05711(.a(new_n4425), .b(new_n257), .O(new_n5905));
  nor2 g05712(.a(new_n5905), .b(new_n4334), .O(new_n5906));
  nor2 g05713(.a(new_n4425), .b(new_n502), .O(new_n5907));
  inv1 g05714(.a(new_n5907), .O(new_n5908));
  nor2 g05715(.a(new_n5908), .b(new_n4732), .O(new_n5909));
  nor2 g05716(.a(new_n5909), .b(new_n5906), .O(new_n5910));
  inv1 g05717(.a(new_n5910), .O(new_n5911));
  nor2 g05718(.a(new_n5911), .b(new_n4099), .O(new_n5912));
  nor2 g05719(.a(new_n5910), .b(new_n4100), .O(new_n5913));
  nor2 g05720(.a(new_n5913), .b(new_n5912), .O(new_n5914));
  nor2 g05721(.a(new_n2660), .b(new_n800), .O(new_n5915));
  inv1 g05722(.a(new_n5915), .O(new_n5916));
  nor2 g05723(.a(new_n2506), .b(new_n847), .O(new_n5917));
  nor2 g05724(.a(new_n2433), .b(new_n941), .O(new_n5918));
  nor2 g05725(.a(new_n5918), .b(new_n5917), .O(new_n5919));
  nor2 g05726(.a(new_n5679), .b(new_n5384), .O(new_n5920));
  nor2 g05727(.a(new_n5920), .b(new_n5919), .O(new_n5921));
  nor2 g05728(.a(new_n5921), .b(new_n5916), .O(new_n5922));
  inv1 g05729(.a(new_n5921), .O(new_n5923));
  nor2 g05730(.a(new_n5923), .b(new_n5915), .O(new_n5924));
  nor2 g05731(.a(new_n5924), .b(new_n5922), .O(new_n5925));
  nor2 g05732(.a(new_n5925), .b(new_n5914), .O(new_n5926));
  inv1 g05733(.a(new_n5914), .O(new_n5927));
  inv1 g05734(.a(new_n5925), .O(new_n5928));
  nor2 g05735(.a(new_n5928), .b(new_n5927), .O(new_n5929));
  nor2 g05736(.a(new_n5929), .b(new_n5926), .O(new_n5930));
  inv1 g05737(.a(new_n5930), .O(new_n5931));
  nor2 g05738(.a(new_n5931), .b(new_n5904), .O(new_n5932));
  nor2 g05739(.a(new_n5930), .b(new_n5903), .O(new_n5933));
  nor2 g05740(.a(new_n5933), .b(new_n5932), .O(new_n5934));
  inv1 g05741(.a(new_n5934), .O(new_n5935));
  nor2 g05742(.a(new_n5935), .b(new_n5886), .O(new_n5936));
  nor2 g05743(.a(new_n5934), .b(new_n5885), .O(new_n5937));
  nor2 g05744(.a(new_n5937), .b(new_n5936), .O(new_n5938));
  inv1 g05745(.a(new_n5938), .O(new_n5939));
  nor2 g05746(.a(new_n5758), .b(new_n5755), .O(new_n5940));
  nor2 g05747(.a(new_n5842), .b(new_n5835), .O(new_n5941));
  nor2 g05748(.a(new_n5941), .b(new_n5940), .O(new_n5942));
  inv1 g05749(.a(new_n5940), .O(new_n5943));
  inv1 g05750(.a(new_n5941), .O(new_n5944));
  nor2 g05751(.a(new_n5944), .b(new_n5943), .O(new_n5945));
  nor2 g05752(.a(new_n5945), .b(new_n5942), .O(new_n5946));
  inv1 g05753(.a(new_n5946), .O(new_n5947));
  nor2 g05754(.a(new_n5947), .b(new_n5939), .O(new_n5948));
  nor2 g05755(.a(new_n5946), .b(new_n5938), .O(new_n5949));
  nor2 g05756(.a(new_n5949), .b(new_n5948), .O(new_n5950));
  nor2 g05757(.a(new_n5950), .b(new_n5866), .O(new_n5951));
  inv1 g05758(.a(new_n5950), .O(new_n5952));
  nor2 g05759(.a(new_n5952), .b(new_n5865), .O(new_n5953));
  nor2 g05760(.a(new_n5953), .b(new_n5951), .O(new_n5954));
  inv1 g05761(.a(new_n5954), .O(new_n5955));
  nor2 g05762(.a(new_n5648), .b(new_n5643), .O(new_n5956));
  inv1 g05763(.a(new_n5956), .O(new_n5957));
  nor2 g05764(.a(new_n5639), .b(new_n5636), .O(new_n5958));
  nor2 g05765(.a(new_n1736), .b(new_n1425), .O(new_n5959));
  nor2 g05766(.a(new_n1647), .b(new_n1493), .O(new_n5960));
  nor2 g05767(.a(new_n5960), .b(new_n5959), .O(new_n5961));
  nor2 g05768(.a(new_n1736), .b(new_n1493), .O(new_n5962));
  inv1 g05769(.a(new_n5962), .O(new_n5963));
  nor2 g05770(.a(new_n5963), .b(new_n5444), .O(new_n5964));
  nor2 g05771(.a(new_n5964), .b(new_n5961), .O(new_n5965));
  nor2 g05772(.a(new_n5965), .b(new_n5432), .O(new_n5966));
  inv1 g05773(.a(new_n5965), .O(new_n5967));
  nor2 g05774(.a(new_n5967), .b(new_n5431), .O(new_n5968));
  nor2 g05775(.a(new_n5968), .b(new_n5966), .O(new_n5969));
  inv1 g05776(.a(new_n5969), .O(new_n5970));
  inv1 g05777(.a(\a[45] ), .O(new_n5971));
  nor2 g05778(.a(new_n5971), .b(new_n198), .O(new_n5972));
  nor2 g05779(.a(new_n5393), .b(new_n196), .O(new_n5973));
  nor2 g05780(.a(new_n4954), .b(new_n214), .O(new_n5974));
  nor2 g05781(.a(new_n5974), .b(new_n5973), .O(new_n5975));
  nor2 g05782(.a(new_n5393), .b(new_n214), .O(new_n5976));
  inv1 g05783(.a(new_n5976), .O(new_n5977));
  nor2 g05784(.a(new_n5977), .b(new_n4959), .O(new_n5978));
  nor2 g05785(.a(new_n5978), .b(new_n5975), .O(new_n5979));
  inv1 g05786(.a(new_n5979), .O(new_n5980));
  nor2 g05787(.a(new_n5980), .b(new_n5972), .O(new_n5981));
  inv1 g05788(.a(new_n5972), .O(new_n5982));
  nor2 g05789(.a(new_n5979), .b(new_n5982), .O(new_n5983));
  nor2 g05790(.a(new_n5983), .b(new_n5981), .O(new_n5984));
  nor2 g05791(.a(new_n4366), .b(new_n295), .O(new_n5985));
  inv1 g05792(.a(new_n5985), .O(new_n5986));
  nor2 g05793(.a(new_n4093), .b(new_n322), .O(new_n5987));
  nor2 g05794(.a(new_n3870), .b(new_n363), .O(new_n5988));
  nor2 g05795(.a(new_n5988), .b(new_n5987), .O(new_n5989));
  nor2 g05796(.a(new_n4093), .b(new_n363), .O(new_n5990));
  inv1 g05797(.a(new_n5990), .O(new_n5991));
  nor2 g05798(.a(new_n5991), .b(new_n5723), .O(new_n5992));
  nor2 g05799(.a(new_n5992), .b(new_n5989), .O(new_n5993));
  nor2 g05800(.a(new_n5993), .b(new_n5986), .O(new_n5994));
  inv1 g05801(.a(new_n5993), .O(new_n5995));
  nor2 g05802(.a(new_n5995), .b(new_n5985), .O(new_n5996));
  nor2 g05803(.a(new_n5996), .b(new_n5994), .O(new_n5997));
  nor2 g05804(.a(new_n5997), .b(new_n5984), .O(new_n5998));
  inv1 g05805(.a(new_n5984), .O(new_n5999));
  inv1 g05806(.a(new_n5997), .O(new_n6000));
  nor2 g05807(.a(new_n6000), .b(new_n5999), .O(new_n6001));
  nor2 g05808(.a(new_n6001), .b(new_n5998), .O(new_n6002));
  nor2 g05809(.a(new_n6002), .b(new_n5970), .O(new_n6003));
  inv1 g05810(.a(new_n6002), .O(new_n6004));
  nor2 g05811(.a(new_n6004), .b(new_n5969), .O(new_n6005));
  nor2 g05812(.a(new_n6005), .b(new_n6003), .O(new_n6006));
  inv1 g05813(.a(new_n6006), .O(new_n6007));
  nor2 g05814(.a(new_n2826), .b(new_n699), .O(new_n6008));
  inv1 g05815(.a(new_n6008), .O(new_n6009));
  nor2 g05816(.a(new_n4682), .b(new_n229), .O(new_n6010));
  nor2 g05817(.a(new_n6010), .b(new_n5713), .O(new_n6011));
  inv1 g05818(.a(new_n6010), .O(new_n6012));
  nor2 g05819(.a(new_n6012), .b(new_n5714), .O(new_n6013));
  nor2 g05820(.a(new_n6013), .b(new_n6011), .O(new_n6014));
  nor2 g05821(.a(new_n6014), .b(new_n6009), .O(new_n6015));
  inv1 g05822(.a(new_n6014), .O(new_n6016));
  nor2 g05823(.a(new_n6016), .b(new_n6008), .O(new_n6017));
  nor2 g05824(.a(new_n6017), .b(new_n6015), .O(new_n6018));
  inv1 g05825(.a(new_n6018), .O(new_n6019));
  nor2 g05826(.a(new_n2184), .b(new_n1086), .O(new_n6020));
  inv1 g05827(.a(new_n6020), .O(new_n6021));
  nor2 g05828(.a(new_n2121), .b(new_n1199), .O(new_n6022));
  nor2 g05829(.a(new_n6022), .b(new_n5691), .O(new_n6023));
  nor2 g05830(.a(new_n2121), .b(new_n1297), .O(new_n6024));
  inv1 g05831(.a(new_n6024), .O(new_n6025));
  nor2 g05832(.a(new_n6025), .b(new_n5371), .O(new_n6026));
  nor2 g05833(.a(new_n6026), .b(new_n6023), .O(new_n6027));
  nor2 g05834(.a(new_n6027), .b(new_n6021), .O(new_n6028));
  inv1 g05835(.a(new_n6027), .O(new_n6029));
  nor2 g05836(.a(new_n6029), .b(new_n6020), .O(new_n6030));
  nor2 g05837(.a(new_n6030), .b(new_n6028), .O(new_n6031));
  nor2 g05838(.a(new_n5730), .b(new_n5725), .O(new_n6032));
  inv1 g05839(.a(new_n6032), .O(new_n6033));
  nor2 g05840(.a(new_n6033), .b(new_n6031), .O(new_n6034));
  inv1 g05841(.a(new_n6031), .O(new_n6035));
  nor2 g05842(.a(new_n6032), .b(new_n6035), .O(new_n6036));
  nor2 g05843(.a(new_n6036), .b(new_n6034), .O(new_n6037));
  nor2 g05844(.a(new_n6037), .b(new_n6019), .O(new_n6038));
  inv1 g05845(.a(new_n6037), .O(new_n6039));
  nor2 g05846(.a(new_n6039), .b(new_n6018), .O(new_n6040));
  nor2 g05847(.a(new_n6040), .b(new_n6038), .O(new_n6041));
  inv1 g05848(.a(new_n6041), .O(new_n6042));
  nor2 g05849(.a(new_n6042), .b(new_n6007), .O(new_n6043));
  nor2 g05850(.a(new_n6041), .b(new_n6006), .O(new_n6044));
  nor2 g05851(.a(new_n6044), .b(new_n6043), .O(new_n6045));
  inv1 g05852(.a(new_n6045), .O(new_n6046));
  nor2 g05853(.a(new_n6046), .b(new_n5958), .O(new_n6047));
  inv1 g05854(.a(new_n5958), .O(new_n6048));
  nor2 g05855(.a(new_n6045), .b(new_n6048), .O(new_n6049));
  nor2 g05856(.a(new_n6049), .b(new_n6047), .O(new_n6050));
  nor2 g05857(.a(new_n6050), .b(new_n5957), .O(new_n6051));
  inv1 g05858(.a(new_n6050), .O(new_n6052));
  nor2 g05859(.a(new_n6052), .b(new_n5956), .O(new_n6053));
  nor2 g05860(.a(new_n6053), .b(new_n6051), .O(new_n6054));
  inv1 g05861(.a(new_n6054), .O(new_n6055));
  nor2 g05862(.a(new_n5628), .b(new_n5622), .O(new_n6056));
  inv1 g05863(.a(new_n6056), .O(new_n6057));
  nor2 g05864(.a(new_n5808), .b(new_n5792), .O(new_n6058));
  inv1 g05865(.a(new_n6058), .O(new_n6059));
  nor2 g05866(.a(new_n6059), .b(new_n6057), .O(new_n6060));
  nor2 g05867(.a(new_n6058), .b(new_n6056), .O(new_n6061));
  nor2 g05868(.a(new_n6061), .b(new_n6060), .O(new_n6062));
  nor2 g05869(.a(new_n5783), .b(new_n5778), .O(new_n6063));
  inv1 g05870(.a(new_n6063), .O(new_n6064));
  nor2 g05871(.a(new_n6064), .b(new_n6062), .O(new_n6065));
  inv1 g05872(.a(new_n6062), .O(new_n6066));
  nor2 g05873(.a(new_n6063), .b(new_n6066), .O(new_n6067));
  nor2 g05874(.a(new_n6067), .b(new_n6065), .O(new_n6068));
  nor2 g05875(.a(new_n5818), .b(new_n5813), .O(new_n6069));
  inv1 g05876(.a(new_n6069), .O(new_n6070));
  nor2 g05877(.a(new_n6070), .b(new_n6068), .O(new_n6071));
  inv1 g05878(.a(new_n6068), .O(new_n6072));
  nor2 g05879(.a(new_n6069), .b(new_n6072), .O(new_n6073));
  nor2 g05880(.a(new_n6073), .b(new_n6071), .O(new_n6074));
  inv1 g05881(.a(new_n6074), .O(new_n6075));
  nor2 g05882(.a(new_n5741), .b(new_n5734), .O(new_n6076));
  nor2 g05883(.a(new_n5671), .b(new_n5664), .O(new_n6077));
  nor2 g05884(.a(new_n6077), .b(new_n6076), .O(new_n6078));
  inv1 g05885(.a(new_n6076), .O(new_n6079));
  inv1 g05886(.a(new_n6077), .O(new_n6080));
  nor2 g05887(.a(new_n6080), .b(new_n6079), .O(new_n6081));
  nor2 g05888(.a(new_n6081), .b(new_n6078), .O(new_n6082));
  nor2 g05889(.a(new_n5719), .b(new_n5712), .O(new_n6083));
  nor2 g05890(.a(new_n6083), .b(new_n6082), .O(new_n6084));
  inv1 g05891(.a(new_n6082), .O(new_n6085));
  inv1 g05892(.a(new_n6083), .O(new_n6086));
  nor2 g05893(.a(new_n6086), .b(new_n6085), .O(new_n6087));
  nor2 g05894(.a(new_n6087), .b(new_n6084), .O(new_n6088));
  inv1 g05895(.a(new_n6088), .O(new_n6089));
  nor2 g05896(.a(new_n5750), .b(new_n5743), .O(new_n6090));
  inv1 g05897(.a(new_n6090), .O(new_n6091));
  nor2 g05898(.a(new_n5706), .b(new_n5699), .O(new_n6092));
  inv1 g05899(.a(new_n6092), .O(new_n6093));
  nor2 g05900(.a(new_n6093), .b(new_n6091), .O(new_n6094));
  nor2 g05901(.a(new_n6092), .b(new_n6090), .O(new_n6095));
  nor2 g05902(.a(new_n6095), .b(new_n6094), .O(new_n6096));
  inv1 g05903(.a(new_n6096), .O(new_n6097));
  nor2 g05904(.a(new_n6097), .b(new_n6089), .O(new_n6098));
  nor2 g05905(.a(new_n6096), .b(new_n6088), .O(new_n6099));
  nor2 g05906(.a(new_n6099), .b(new_n6098), .O(new_n6100));
  inv1 g05907(.a(new_n6100), .O(new_n6101));
  nor2 g05908(.a(new_n6101), .b(new_n6075), .O(new_n6102));
  nor2 g05909(.a(new_n6100), .b(new_n6074), .O(new_n6103));
  nor2 g05910(.a(new_n6103), .b(new_n6102), .O(new_n6104));
  inv1 g05911(.a(new_n6104), .O(new_n6105));
  nor2 g05912(.a(new_n6105), .b(new_n6055), .O(new_n6106));
  nor2 g05913(.a(new_n6104), .b(new_n6054), .O(new_n6107));
  nor2 g05914(.a(new_n6107), .b(new_n6106), .O(new_n6108));
  inv1 g05915(.a(new_n6108), .O(new_n6109));
  nor2 g05916(.a(new_n6109), .b(new_n5955), .O(new_n6110));
  nor2 g05917(.a(new_n6108), .b(new_n5954), .O(new_n6111));
  nor2 g05918(.a(new_n6111), .b(new_n6110), .O(new_n6112));
  inv1 g05919(.a(new_n6112), .O(new_n6113));
  nor2 g05920(.a(new_n6113), .b(new_n5864), .O(new_n6114));
  inv1 g05921(.a(new_n5864), .O(new_n6115));
  nor2 g05922(.a(new_n6112), .b(new_n6115), .O(new_n6116));
  nor2 g05923(.a(new_n6116), .b(new_n6114), .O(new_n6117));
  inv1 g05924(.a(new_n6117), .O(new_n6118));
  nor2 g05925(.a(new_n5859), .b(new_n5855), .O(new_n6119));
  nor2 g05926(.a(new_n6119), .b(new_n6118), .O(new_n6120));
  inv1 g05927(.a(new_n6119), .O(new_n6121));
  nor2 g05928(.a(new_n6121), .b(new_n6117), .O(new_n6122));
  nor2 g05929(.a(new_n6122), .b(new_n6120), .O(new_n6123));
  inv1 g05930(.a(new_n6123), .O(\asquared[46] ));
  nor2 g05931(.a(new_n6110), .b(new_n5953), .O(new_n6125));
  inv1 g05932(.a(new_n6125), .O(new_n6126));
  nor2 g05933(.a(new_n6106), .b(new_n6053), .O(new_n6127));
  nor2 g05934(.a(new_n6102), .b(new_n6073), .O(new_n6128));
  inv1 g05935(.a(new_n6128), .O(new_n6129));
  nor2 g05936(.a(new_n6047), .b(new_n6043), .O(new_n6130));
  inv1 g05937(.a(new_n6130), .O(new_n6131));
  nor2 g05938(.a(new_n6131), .b(new_n6129), .O(new_n6132));
  nor2 g05939(.a(new_n6130), .b(new_n6128), .O(new_n6133));
  nor2 g05940(.a(new_n6133), .b(new_n6132), .O(new_n6134));
  inv1 g05941(.a(new_n6134), .O(new_n6135));
  nor2 g05942(.a(new_n6087), .b(new_n6081), .O(new_n6136));
  inv1 g05943(.a(new_n6136), .O(new_n6137));
  nor2 g05944(.a(new_n2826), .b(new_n800), .O(new_n6138));
  nor2 g05945(.a(new_n4954), .b(new_n229), .O(new_n6139));
  nor2 g05946(.a(new_n6139), .b(new_n6138), .O(new_n6140));
  inv1 g05947(.a(new_n3945), .O(new_n6141));
  nor2 g05948(.a(new_n4954), .b(new_n800), .O(new_n6142));
  inv1 g05949(.a(new_n6142), .O(new_n6143));
  nor2 g05950(.a(new_n6143), .b(new_n6141), .O(new_n6144));
  nor2 g05951(.a(new_n6144), .b(new_n6140), .O(new_n6145));
  inv1 g05952(.a(new_n6145), .O(new_n6146));
  nor2 g05953(.a(new_n6146), .b(new_n5800), .O(new_n6147));
  nor2 g05954(.a(new_n6145), .b(new_n5801), .O(new_n6148));
  nor2 g05955(.a(new_n6148), .b(new_n6147), .O(new_n6149));
  nor2 g05956(.a(new_n3057), .b(new_n699), .O(new_n6150));
  inv1 g05957(.a(new_n6150), .O(new_n6151));
  nor2 g05958(.a(new_n4682), .b(new_n257), .O(new_n6152));
  nor2 g05959(.a(new_n3231), .b(new_n613), .O(new_n6153));
  nor2 g05960(.a(new_n6153), .b(new_n6152), .O(new_n6154));
  inv1 g05961(.a(new_n6152), .O(new_n6155));
  inv1 g05962(.a(new_n6153), .O(new_n6156));
  nor2 g05963(.a(new_n6156), .b(new_n6155), .O(new_n6157));
  nor2 g05964(.a(new_n6157), .b(new_n6154), .O(new_n6158));
  nor2 g05965(.a(new_n6158), .b(new_n6151), .O(new_n6159));
  inv1 g05966(.a(new_n6158), .O(new_n6160));
  nor2 g05967(.a(new_n6160), .b(new_n6150), .O(new_n6161));
  nor2 g05968(.a(new_n6161), .b(new_n6159), .O(new_n6162));
  nor2 g05969(.a(new_n6162), .b(new_n6149), .O(new_n6163));
  inv1 g05970(.a(new_n6149), .O(new_n6164));
  inv1 g05971(.a(new_n6162), .O(new_n6165));
  nor2 g05972(.a(new_n6165), .b(new_n6164), .O(new_n6166));
  nor2 g05973(.a(new_n6166), .b(new_n6163), .O(new_n6167));
  nor2 g05974(.a(new_n6167), .b(new_n6137), .O(new_n6168));
  inv1 g05975(.a(new_n6167), .O(new_n6169));
  nor2 g05976(.a(new_n6169), .b(new_n6136), .O(new_n6170));
  nor2 g05977(.a(new_n6170), .b(new_n6168), .O(new_n6171));
  inv1 g05978(.a(new_n6171), .O(new_n6172));
  nor2 g05979(.a(new_n5924), .b(new_n5919), .O(new_n6173));
  nor2 g05980(.a(new_n6030), .b(new_n6023), .O(new_n6174));
  nor2 g05981(.a(new_n6174), .b(new_n6173), .O(new_n6175));
  inv1 g05982(.a(new_n6173), .O(new_n6176));
  inv1 g05983(.a(new_n6174), .O(new_n6177));
  nor2 g05984(.a(new_n6177), .b(new_n6176), .O(new_n6178));
  nor2 g05985(.a(new_n6178), .b(new_n6175), .O(new_n6179));
  nor2 g05986(.a(new_n5912), .b(new_n5906), .O(new_n6180));
  nor2 g05987(.a(new_n6180), .b(new_n6179), .O(new_n6181));
  inv1 g05988(.a(new_n6179), .O(new_n6182));
  inv1 g05989(.a(new_n6180), .O(new_n6183));
  nor2 g05990(.a(new_n6183), .b(new_n6182), .O(new_n6184));
  nor2 g05991(.a(new_n6184), .b(new_n6181), .O(new_n6185));
  nor2 g05992(.a(new_n6067), .b(new_n6061), .O(new_n6186));
  inv1 g05993(.a(new_n6186), .O(new_n6187));
  nor2 g05994(.a(new_n6187), .b(new_n6185), .O(new_n6188));
  inv1 g05995(.a(new_n6185), .O(new_n6189));
  nor2 g05996(.a(new_n6186), .b(new_n6189), .O(new_n6190));
  nor2 g05997(.a(new_n6190), .b(new_n6188), .O(new_n6191));
  inv1 g05998(.a(new_n6191), .O(new_n6192));
  nor2 g05999(.a(new_n6192), .b(new_n6172), .O(new_n6193));
  nor2 g06000(.a(new_n6191), .b(new_n6171), .O(new_n6194));
  nor2 g06001(.a(new_n6194), .b(new_n6193), .O(new_n6195));
  inv1 g06002(.a(new_n6195), .O(new_n6196));
  nor2 g06003(.a(new_n6196), .b(new_n6135), .O(new_n6197));
  nor2 g06004(.a(new_n6195), .b(new_n6134), .O(new_n6198));
  nor2 g06005(.a(new_n6198), .b(new_n6197), .O(new_n6199));
  inv1 g06006(.a(new_n6199), .O(new_n6200));
  nor2 g06007(.a(new_n6200), .b(new_n6127), .O(new_n6201));
  inv1 g06008(.a(new_n6127), .O(new_n6202));
  nor2 g06009(.a(new_n6199), .b(new_n6202), .O(new_n6203));
  nor2 g06010(.a(new_n6203), .b(new_n6201), .O(new_n6204));
  nor2 g06011(.a(new_n6204), .b(new_n6126), .O(new_n6205));
  inv1 g06012(.a(new_n6204), .O(new_n6206));
  nor2 g06013(.a(new_n6206), .b(new_n6125), .O(new_n6207));
  nor2 g06014(.a(new_n6207), .b(new_n6205), .O(new_n6208));
  nor2 g06015(.a(new_n5948), .b(new_n5942), .O(new_n6209));
  nor2 g06016(.a(new_n6098), .b(new_n6095), .O(new_n6210));
  nor2 g06017(.a(new_n3533), .b(new_n569), .O(new_n6211));
  inv1 g06018(.a(new_n6211), .O(new_n6212));
  nor2 g06019(.a(new_n4425), .b(new_n295), .O(new_n6213));
  nor2 g06020(.a(new_n4366), .b(new_n322), .O(new_n6214));
  nor2 g06021(.a(new_n6214), .b(new_n6213), .O(new_n6215));
  nor2 g06022(.a(new_n4425), .b(new_n322), .O(new_n6216));
  inv1 g06023(.a(new_n6216), .O(new_n6217));
  nor2 g06024(.a(new_n6217), .b(new_n5986), .O(new_n6218));
  nor2 g06025(.a(new_n6218), .b(new_n6215), .O(new_n6219));
  nor2 g06026(.a(new_n6219), .b(new_n6212), .O(new_n6220));
  inv1 g06027(.a(new_n6219), .O(new_n6221));
  nor2 g06028(.a(new_n6221), .b(new_n6211), .O(new_n6222));
  nor2 g06029(.a(new_n6222), .b(new_n6220), .O(new_n6223));
  nor2 g06030(.a(new_n5900), .b(new_n5891), .O(new_n6224));
  nor2 g06031(.a(new_n2660), .b(new_n847), .O(new_n6225));
  inv1 g06032(.a(new_n6225), .O(new_n6226));
  nor2 g06033(.a(new_n2433), .b(new_n1086), .O(new_n6227));
  nor2 g06034(.a(new_n6227), .b(new_n5678), .O(new_n6228));
  inv1 g06035(.a(new_n5918), .O(new_n6229));
  nor2 g06036(.a(new_n2506), .b(new_n1086), .O(new_n6230));
  inv1 g06037(.a(new_n6230), .O(new_n6231));
  nor2 g06038(.a(new_n6231), .b(new_n6229), .O(new_n6232));
  nor2 g06039(.a(new_n6232), .b(new_n6228), .O(new_n6233));
  nor2 g06040(.a(new_n6233), .b(new_n6226), .O(new_n6234));
  inv1 g06041(.a(new_n6233), .O(new_n6235));
  nor2 g06042(.a(new_n6235), .b(new_n6225), .O(new_n6236));
  nor2 g06043(.a(new_n6236), .b(new_n6234), .O(new_n6237));
  nor2 g06044(.a(new_n6237), .b(new_n6224), .O(new_n6238));
  inv1 g06045(.a(new_n6224), .O(new_n6239));
  inv1 g06046(.a(new_n6237), .O(new_n6240));
  nor2 g06047(.a(new_n6240), .b(new_n6239), .O(new_n6241));
  nor2 g06048(.a(new_n6241), .b(new_n6238), .O(new_n6242));
  inv1 g06049(.a(new_n6242), .O(new_n6243));
  nor2 g06050(.a(new_n6243), .b(new_n6223), .O(new_n6244));
  inv1 g06051(.a(new_n6223), .O(new_n6245));
  nor2 g06052(.a(new_n6242), .b(new_n6245), .O(new_n6246));
  nor2 g06053(.a(new_n6246), .b(new_n6244), .O(new_n6247));
  inv1 g06054(.a(new_n6247), .O(new_n6248));
  nor2 g06055(.a(new_n2184), .b(new_n1199), .O(new_n6249));
  inv1 g06056(.a(new_n6249), .O(new_n6250));
  nor2 g06057(.a(new_n1903), .b(new_n1425), .O(new_n6251));
  nor2 g06058(.a(new_n6251), .b(new_n6024), .O(new_n6252));
  nor2 g06059(.a(new_n2121), .b(new_n1425), .O(new_n6253));
  inv1 g06060(.a(new_n6253), .O(new_n6254));
  nor2 g06061(.a(new_n6254), .b(new_n5692), .O(new_n6255));
  nor2 g06062(.a(new_n6255), .b(new_n6252), .O(new_n6256));
  nor2 g06063(.a(new_n6256), .b(new_n6250), .O(new_n6257));
  inv1 g06064(.a(new_n6256), .O(new_n6258));
  nor2 g06065(.a(new_n6258), .b(new_n6249), .O(new_n6259));
  nor2 g06066(.a(new_n6259), .b(new_n6257), .O(new_n6260));
  inv1 g06067(.a(new_n6260), .O(new_n6261));
  nor2 g06068(.a(new_n3870), .b(new_n438), .O(new_n6262));
  nor2 g06069(.a(new_n6262), .b(new_n5008), .O(new_n6263));
  nor2 g06070(.a(new_n3870), .b(new_n502), .O(new_n6264));
  inv1 g06071(.a(new_n6264), .O(new_n6265));
  nor2 g06072(.a(new_n6265), .b(new_n5432), .O(new_n6266));
  nor2 g06073(.a(new_n6266), .b(new_n6263), .O(new_n6267));
  nor2 g06074(.a(new_n6267), .b(new_n5991), .O(new_n6268));
  inv1 g06075(.a(new_n6267), .O(new_n6269));
  nor2 g06076(.a(new_n6269), .b(new_n5990), .O(new_n6270));
  nor2 g06077(.a(new_n6270), .b(new_n6268), .O(new_n6271));
  nor2 g06078(.a(new_n5393), .b(new_n203), .O(new_n6272));
  inv1 g06079(.a(new_n6272), .O(new_n6273));
  inv1 g06080(.a(\a[46] ), .O(new_n6274));
  nor2 g06081(.a(new_n6274), .b(new_n198), .O(new_n6275));
  nor2 g06082(.a(new_n5178), .b(new_n214), .O(new_n6276));
  nor2 g06083(.a(new_n6276), .b(new_n6275), .O(new_n6277));
  inv1 g06084(.a(new_n6275), .O(new_n6278));
  inv1 g06085(.a(new_n6276), .O(new_n6279));
  nor2 g06086(.a(new_n6279), .b(new_n6278), .O(new_n6280));
  nor2 g06087(.a(new_n6280), .b(new_n6277), .O(new_n6281));
  nor2 g06088(.a(new_n6281), .b(new_n6273), .O(new_n6282));
  inv1 g06089(.a(new_n6281), .O(new_n6283));
  nor2 g06090(.a(new_n6283), .b(new_n6272), .O(new_n6284));
  nor2 g06091(.a(new_n6284), .b(new_n6282), .O(new_n6285));
  nor2 g06092(.a(new_n6285), .b(new_n6271), .O(new_n6286));
  inv1 g06093(.a(new_n6271), .O(new_n6287));
  inv1 g06094(.a(new_n6285), .O(new_n6288));
  nor2 g06095(.a(new_n6288), .b(new_n6287), .O(new_n6289));
  nor2 g06096(.a(new_n6289), .b(new_n6286), .O(new_n6290));
  nor2 g06097(.a(new_n6290), .b(new_n6261), .O(new_n6291));
  inv1 g06098(.a(new_n6290), .O(new_n6292));
  nor2 g06099(.a(new_n6292), .b(new_n6260), .O(new_n6293));
  nor2 g06100(.a(new_n6293), .b(new_n6291), .O(new_n6294));
  inv1 g06101(.a(new_n6294), .O(new_n6295));
  nor2 g06102(.a(new_n6295), .b(new_n6248), .O(new_n6296));
  nor2 g06103(.a(new_n6294), .b(new_n6247), .O(new_n6297));
  nor2 g06104(.a(new_n6297), .b(new_n6296), .O(new_n6298));
  inv1 g06105(.a(new_n6298), .O(new_n6299));
  nor2 g06106(.a(new_n6299), .b(new_n6210), .O(new_n6300));
  inv1 g06107(.a(new_n6210), .O(new_n6301));
  nor2 g06108(.a(new_n6298), .b(new_n6301), .O(new_n6302));
  nor2 g06109(.a(new_n6302), .b(new_n6300), .O(new_n6303));
  inv1 g06110(.a(new_n6303), .O(new_n6304));
  nor2 g06111(.a(new_n6304), .b(new_n6209), .O(new_n6305));
  inv1 g06112(.a(new_n6209), .O(new_n6306));
  nor2 g06113(.a(new_n6303), .b(new_n6306), .O(new_n6307));
  nor2 g06114(.a(new_n6307), .b(new_n6305), .O(new_n6308));
  inv1 g06115(.a(new_n6308), .O(new_n6309));
  nor2 g06116(.a(new_n6005), .b(new_n5998), .O(new_n6310));
  inv1 g06117(.a(new_n6310), .O(new_n6311));
  nor2 g06118(.a(new_n6040), .b(new_n6034), .O(new_n6312));
  inv1 g06119(.a(new_n6312), .O(new_n6313));
  nor2 g06120(.a(new_n6313), .b(new_n6311), .O(new_n6314));
  nor2 g06121(.a(new_n6312), .b(new_n6310), .O(new_n6315));
  nor2 g06122(.a(new_n6315), .b(new_n6314), .O(new_n6316));
  nor2 g06123(.a(new_n5932), .b(new_n5926), .O(new_n6317));
  inv1 g06124(.a(new_n6317), .O(new_n6318));
  nor2 g06125(.a(new_n6318), .b(new_n6316), .O(new_n6319));
  inv1 g06126(.a(new_n6316), .O(new_n6320));
  nor2 g06127(.a(new_n6317), .b(new_n6320), .O(new_n6321));
  nor2 g06128(.a(new_n6321), .b(new_n6319), .O(new_n6322));
  inv1 g06129(.a(new_n6322), .O(new_n6323));
  nor2 g06130(.a(new_n5936), .b(new_n5884), .O(new_n6324));
  nor2 g06131(.a(new_n6017), .b(new_n6011), .O(new_n6325));
  nor2 g06132(.a(new_n5981), .b(new_n5975), .O(new_n6326));
  nor2 g06133(.a(new_n6326), .b(new_n6325), .O(new_n6327));
  inv1 g06134(.a(new_n6325), .O(new_n6328));
  inv1 g06135(.a(new_n6326), .O(new_n6329));
  nor2 g06136(.a(new_n6329), .b(new_n6328), .O(new_n6330));
  nor2 g06137(.a(new_n6330), .b(new_n6327), .O(new_n6331));
  nor2 g06138(.a(new_n5996), .b(new_n5989), .O(new_n6332));
  nor2 g06139(.a(new_n6332), .b(new_n6331), .O(new_n6333));
  inv1 g06140(.a(new_n6331), .O(new_n6334));
  inv1 g06141(.a(new_n6332), .O(new_n6335));
  nor2 g06142(.a(new_n6335), .b(new_n6334), .O(new_n6336));
  nor2 g06143(.a(new_n6336), .b(new_n6333), .O(new_n6337));
  inv1 g06144(.a(new_n6337), .O(new_n6338));
  nor2 g06145(.a(new_n5878), .b(new_n5872), .O(new_n6339));
  inv1 g06146(.a(new_n5894), .O(new_n6340));
  nor2 g06147(.a(new_n5971), .b(new_n194), .O(new_n6341));
  nor2 g06148(.a(new_n6341), .b(new_n5962), .O(new_n6342));
  inv1 g06149(.a(new_n6341), .O(new_n6343));
  nor2 g06150(.a(new_n6343), .b(new_n5963), .O(new_n6344));
  nor2 g06151(.a(new_n6344), .b(new_n6342), .O(new_n6345));
  inv1 g06152(.a(new_n6345), .O(new_n6346));
  nor2 g06153(.a(new_n6346), .b(new_n6340), .O(new_n6347));
  nor2 g06154(.a(new_n6345), .b(new_n5894), .O(new_n6348));
  nor2 g06155(.a(new_n6348), .b(new_n6347), .O(new_n6349));
  inv1 g06156(.a(new_n6349), .O(new_n6350));
  nor2 g06157(.a(new_n5968), .b(new_n5961), .O(new_n6351));
  inv1 g06158(.a(new_n6351), .O(new_n6352));
  nor2 g06159(.a(new_n6352), .b(new_n6350), .O(new_n6353));
  nor2 g06160(.a(new_n6351), .b(new_n6349), .O(new_n6354));
  nor2 g06161(.a(new_n6354), .b(new_n6353), .O(new_n6355));
  inv1 g06162(.a(new_n6355), .O(new_n6356));
  nor2 g06163(.a(new_n6356), .b(new_n6339), .O(new_n6357));
  inv1 g06164(.a(new_n6339), .O(new_n6358));
  nor2 g06165(.a(new_n6355), .b(new_n6358), .O(new_n6359));
  nor2 g06166(.a(new_n6359), .b(new_n6357), .O(new_n6360));
  inv1 g06167(.a(new_n6360), .O(new_n6361));
  nor2 g06168(.a(new_n6361), .b(new_n6338), .O(new_n6362));
  nor2 g06169(.a(new_n6360), .b(new_n6337), .O(new_n6363));
  nor2 g06170(.a(new_n6363), .b(new_n6362), .O(new_n6364));
  inv1 g06171(.a(new_n6364), .O(new_n6365));
  nor2 g06172(.a(new_n6365), .b(new_n6324), .O(new_n6366));
  inv1 g06173(.a(new_n6324), .O(new_n6367));
  nor2 g06174(.a(new_n6364), .b(new_n6367), .O(new_n6368));
  nor2 g06175(.a(new_n6368), .b(new_n6366), .O(new_n6369));
  inv1 g06176(.a(new_n6369), .O(new_n6370));
  nor2 g06177(.a(new_n6370), .b(new_n6323), .O(new_n6371));
  nor2 g06178(.a(new_n6369), .b(new_n6322), .O(new_n6372));
  nor2 g06179(.a(new_n6372), .b(new_n6371), .O(new_n6373));
  inv1 g06180(.a(new_n6373), .O(new_n6374));
  nor2 g06181(.a(new_n6374), .b(new_n6309), .O(new_n6375));
  nor2 g06182(.a(new_n6373), .b(new_n6308), .O(new_n6376));
  nor2 g06183(.a(new_n6376), .b(new_n6375), .O(new_n6377));
  nor2 g06184(.a(new_n6377), .b(new_n6208), .O(new_n6378));
  inv1 g06185(.a(new_n6208), .O(new_n6379));
  inv1 g06186(.a(new_n6377), .O(new_n6380));
  nor2 g06187(.a(new_n6380), .b(new_n6379), .O(new_n6381));
  nor2 g06188(.a(new_n6381), .b(new_n6378), .O(new_n6382));
  inv1 g06189(.a(new_n6382), .O(new_n6383));
  nor2 g06190(.a(new_n6120), .b(new_n6116), .O(new_n6384));
  nor2 g06191(.a(new_n6384), .b(new_n6383), .O(new_n6385));
  inv1 g06192(.a(new_n6384), .O(new_n6386));
  nor2 g06193(.a(new_n6386), .b(new_n6382), .O(new_n6387));
  nor2 g06194(.a(new_n6387), .b(new_n6385), .O(new_n6388));
  inv1 g06195(.a(new_n6388), .O(\asquared[47] ));
  nor2 g06196(.a(new_n6207), .b(new_n6201), .O(new_n6390));
  nor2 g06197(.a(new_n6197), .b(new_n6133), .O(new_n6391));
  inv1 g06198(.a(new_n6391), .O(new_n6392));
  nor2 g06199(.a(new_n6371), .b(new_n6366), .O(new_n6393));
  inv1 g06200(.a(new_n6393), .O(new_n6394));
  nor2 g06201(.a(new_n6394), .b(new_n6392), .O(new_n6395));
  nor2 g06202(.a(new_n6393), .b(new_n6391), .O(new_n6396));
  nor2 g06203(.a(new_n6396), .b(new_n6395), .O(new_n6397));
  inv1 g06204(.a(new_n6397), .O(new_n6398));
  nor2 g06205(.a(new_n6259), .b(new_n6252), .O(new_n6399));
  nor2 g06206(.a(new_n6147), .b(new_n6140), .O(new_n6400));
  nor2 g06207(.a(new_n6400), .b(new_n6399), .O(new_n6401));
  inv1 g06208(.a(new_n6399), .O(new_n6402));
  inv1 g06209(.a(new_n6400), .O(new_n6403));
  nor2 g06210(.a(new_n6403), .b(new_n6402), .O(new_n6404));
  nor2 g06211(.a(new_n6404), .b(new_n6401), .O(new_n6405));
  nor2 g06212(.a(new_n6284), .b(new_n6277), .O(new_n6406));
  nor2 g06213(.a(new_n6406), .b(new_n6405), .O(new_n6407));
  inv1 g06214(.a(new_n6405), .O(new_n6408));
  inv1 g06215(.a(new_n6406), .O(new_n6409));
  nor2 g06216(.a(new_n6409), .b(new_n6408), .O(new_n6410));
  nor2 g06217(.a(new_n6410), .b(new_n6407), .O(new_n6411));
  nor2 g06218(.a(new_n6293), .b(new_n6286), .O(new_n6412));
  inv1 g06219(.a(new_n6412), .O(new_n6413));
  nor2 g06220(.a(new_n6413), .b(new_n6411), .O(new_n6414));
  inv1 g06221(.a(new_n6411), .O(new_n6415));
  nor2 g06222(.a(new_n6412), .b(new_n6415), .O(new_n6416));
  nor2 g06223(.a(new_n6416), .b(new_n6414), .O(new_n6417));
  nor2 g06224(.a(new_n6170), .b(new_n6163), .O(new_n6418));
  inv1 g06225(.a(new_n6418), .O(new_n6419));
  nor2 g06226(.a(new_n6419), .b(new_n6417), .O(new_n6420));
  inv1 g06227(.a(new_n6417), .O(new_n6421));
  nor2 g06228(.a(new_n6418), .b(new_n6421), .O(new_n6422));
  nor2 g06229(.a(new_n6422), .b(new_n6420), .O(new_n6423));
  inv1 g06230(.a(new_n6423), .O(new_n6424));
  nor2 g06231(.a(new_n6300), .b(new_n6296), .O(new_n6425));
  nor2 g06232(.a(new_n6193), .b(new_n6190), .O(new_n6426));
  nor2 g06233(.a(new_n6426), .b(new_n6425), .O(new_n6427));
  inv1 g06234(.a(new_n6425), .O(new_n6428));
  inv1 g06235(.a(new_n6426), .O(new_n6429));
  nor2 g06236(.a(new_n6429), .b(new_n6428), .O(new_n6430));
  nor2 g06237(.a(new_n6430), .b(new_n6427), .O(new_n6431));
  inv1 g06238(.a(new_n6431), .O(new_n6432));
  nor2 g06239(.a(new_n6432), .b(new_n6424), .O(new_n6433));
  nor2 g06240(.a(new_n6431), .b(new_n6423), .O(new_n6434));
  nor2 g06241(.a(new_n6434), .b(new_n6433), .O(new_n6435));
  inv1 g06242(.a(new_n6435), .O(new_n6436));
  nor2 g06243(.a(new_n6436), .b(new_n6398), .O(new_n6437));
  nor2 g06244(.a(new_n6435), .b(new_n6397), .O(new_n6438));
  nor2 g06245(.a(new_n6438), .b(new_n6437), .O(new_n6439));
  inv1 g06246(.a(new_n6439), .O(new_n6440));
  nor2 g06247(.a(new_n6375), .b(new_n6305), .O(new_n6441));
  nor2 g06248(.a(new_n6184), .b(new_n6178), .O(new_n6442));
  inv1 g06249(.a(new_n6442), .O(new_n6443));
  nor2 g06250(.a(new_n6353), .b(new_n6347), .O(new_n6444));
  nor2 g06251(.a(new_n3533), .b(new_n613), .O(new_n6445));
  inv1 g06252(.a(new_n6445), .O(new_n6446));
  nor2 g06253(.a(new_n3722), .b(new_n569), .O(new_n6447));
  nor2 g06254(.a(new_n4682), .b(new_n295), .O(new_n6448));
  nor2 g06255(.a(new_n6448), .b(new_n6447), .O(new_n6449));
  nor2 g06256(.a(new_n4682), .b(new_n569), .O(new_n6450));
  inv1 g06257(.a(new_n6450), .O(new_n6451));
  nor2 g06258(.a(new_n6451), .b(new_n5263), .O(new_n6452));
  nor2 g06259(.a(new_n6452), .b(new_n6449), .O(new_n6453));
  nor2 g06260(.a(new_n6453), .b(new_n6446), .O(new_n6454));
  inv1 g06261(.a(new_n6453), .O(new_n6455));
  nor2 g06262(.a(new_n6455), .b(new_n6445), .O(new_n6456));
  nor2 g06263(.a(new_n6456), .b(new_n6454), .O(new_n6457));
  nor2 g06264(.a(new_n6457), .b(new_n6444), .O(new_n6458));
  inv1 g06265(.a(new_n6444), .O(new_n6459));
  inv1 g06266(.a(new_n6457), .O(new_n6460));
  nor2 g06267(.a(new_n6460), .b(new_n6459), .O(new_n6461));
  nor2 g06268(.a(new_n6461), .b(new_n6458), .O(new_n6462));
  nor2 g06269(.a(new_n6462), .b(new_n6443), .O(new_n6463));
  inv1 g06270(.a(new_n6462), .O(new_n6464));
  nor2 g06271(.a(new_n6464), .b(new_n6442), .O(new_n6465));
  nor2 g06272(.a(new_n6465), .b(new_n6463), .O(new_n6466));
  nor2 g06273(.a(new_n6362), .b(new_n6357), .O(new_n6467));
  inv1 g06274(.a(new_n6467), .O(new_n6468));
  nor2 g06275(.a(new_n6468), .b(new_n6466), .O(new_n6469));
  inv1 g06276(.a(new_n6466), .O(new_n6470));
  nor2 g06277(.a(new_n6467), .b(new_n6470), .O(new_n6471));
  nor2 g06278(.a(new_n6471), .b(new_n6469), .O(new_n6472));
  nor2 g06279(.a(new_n6321), .b(new_n6315), .O(new_n6473));
  inv1 g06280(.a(new_n6473), .O(new_n6474));
  nor2 g06281(.a(new_n6474), .b(new_n6472), .O(new_n6475));
  inv1 g06282(.a(new_n6472), .O(new_n6476));
  nor2 g06283(.a(new_n6473), .b(new_n6476), .O(new_n6477));
  nor2 g06284(.a(new_n6477), .b(new_n6475), .O(new_n6478));
  inv1 g06285(.a(new_n6478), .O(new_n6479));
  nor2 g06286(.a(new_n6161), .b(new_n6154), .O(new_n6480));
  nor2 g06287(.a(new_n6236), .b(new_n6228), .O(new_n6481));
  nor2 g06288(.a(new_n6481), .b(new_n6480), .O(new_n6482));
  inv1 g06289(.a(new_n6480), .O(new_n6483));
  inv1 g06290(.a(new_n6481), .O(new_n6484));
  nor2 g06291(.a(new_n6484), .b(new_n6483), .O(new_n6485));
  nor2 g06292(.a(new_n6485), .b(new_n6482), .O(new_n6486));
  inv1 g06293(.a(new_n6486), .O(new_n6487));
  nor2 g06294(.a(new_n5796), .b(new_n203), .O(new_n6488));
  inv1 g06295(.a(new_n6488), .O(new_n6489));
  nor2 g06296(.a(new_n3057), .b(new_n800), .O(new_n6490));
  nor2 g06297(.a(new_n6490), .b(new_n5976), .O(new_n6491));
  nor2 g06298(.a(new_n5393), .b(new_n800), .O(new_n6492));
  inv1 g06299(.a(new_n6492), .O(new_n6493));
  nor2 g06300(.a(new_n6493), .b(new_n3899), .O(new_n6494));
  nor2 g06301(.a(new_n6494), .b(new_n6491), .O(new_n6495));
  nor2 g06302(.a(new_n6495), .b(new_n6489), .O(new_n6496));
  inv1 g06303(.a(new_n6495), .O(new_n6497));
  nor2 g06304(.a(new_n6497), .b(new_n6488), .O(new_n6498));
  nor2 g06305(.a(new_n6498), .b(new_n6496), .O(new_n6499));
  nor2 g06306(.a(new_n6499), .b(new_n6487), .O(new_n6500));
  inv1 g06307(.a(new_n6499), .O(new_n6501));
  nor2 g06308(.a(new_n6501), .b(new_n6486), .O(new_n6502));
  nor2 g06309(.a(new_n6502), .b(new_n6500), .O(new_n6503));
  inv1 g06310(.a(new_n6503), .O(new_n6504));
  nor2 g06311(.a(new_n5178), .b(new_n229), .O(new_n6505));
  inv1 g06312(.a(new_n6505), .O(new_n6506));
  nor2 g06313(.a(new_n4954), .b(new_n257), .O(new_n6507));
  nor2 g06314(.a(new_n3231), .b(new_n699), .O(new_n6508));
  nor2 g06315(.a(new_n6508), .b(new_n6507), .O(new_n6509));
  nor2 g06316(.a(new_n4954), .b(new_n699), .O(new_n6510));
  inv1 g06317(.a(new_n6510), .O(new_n6511));
  nor2 g06318(.a(new_n6511), .b(new_n4525), .O(new_n6512));
  nor2 g06319(.a(new_n6512), .b(new_n6509), .O(new_n6513));
  nor2 g06320(.a(new_n6513), .b(new_n6506), .O(new_n6514));
  inv1 g06321(.a(new_n6513), .O(new_n6515));
  nor2 g06322(.a(new_n6515), .b(new_n6505), .O(new_n6516));
  nor2 g06323(.a(new_n6516), .b(new_n6514), .O(new_n6517));
  inv1 g06324(.a(new_n6517), .O(new_n6518));
  nor2 g06325(.a(new_n4366), .b(new_n363), .O(new_n6519));
  nor2 g06326(.a(new_n6519), .b(new_n6264), .O(new_n6520));
  inv1 g06327(.a(new_n5988), .O(new_n6521));
  nor2 g06328(.a(new_n4366), .b(new_n502), .O(new_n6522));
  inv1 g06329(.a(new_n6522), .O(new_n6523));
  nor2 g06330(.a(new_n6523), .b(new_n6521), .O(new_n6524));
  nor2 g06331(.a(new_n6524), .b(new_n6520), .O(new_n6525));
  inv1 g06332(.a(new_n6525), .O(new_n6526));
  nor2 g06333(.a(new_n6526), .b(new_n6216), .O(new_n6527));
  nor2 g06334(.a(new_n6525), .b(new_n6217), .O(new_n6528));
  nor2 g06335(.a(new_n6528), .b(new_n6527), .O(new_n6529));
  nor2 g06336(.a(new_n4093), .b(new_n438), .O(new_n6530));
  inv1 g06337(.a(new_n6530), .O(new_n6531));
  nor2 g06338(.a(new_n1736), .b(new_n1647), .O(new_n6532));
  nor2 g06339(.a(new_n1903), .b(new_n1493), .O(new_n6533));
  nor2 g06340(.a(new_n6533), .b(new_n6532), .O(new_n6534));
  nor2 g06341(.a(new_n1903), .b(new_n1647), .O(new_n6535));
  inv1 g06342(.a(new_n6535), .O(new_n6536));
  nor2 g06343(.a(new_n6536), .b(new_n5963), .O(new_n6537));
  nor2 g06344(.a(new_n6537), .b(new_n6534), .O(new_n6538));
  nor2 g06345(.a(new_n6538), .b(new_n6531), .O(new_n6539));
  inv1 g06346(.a(new_n6538), .O(new_n6540));
  nor2 g06347(.a(new_n6540), .b(new_n6530), .O(new_n6541));
  nor2 g06348(.a(new_n6541), .b(new_n6539), .O(new_n6542));
  nor2 g06349(.a(new_n6542), .b(new_n6529), .O(new_n6543));
  inv1 g06350(.a(new_n6529), .O(new_n6544));
  inv1 g06351(.a(new_n6542), .O(new_n6545));
  nor2 g06352(.a(new_n6545), .b(new_n6544), .O(new_n6546));
  nor2 g06353(.a(new_n6546), .b(new_n6543), .O(new_n6547));
  nor2 g06354(.a(new_n6547), .b(new_n6518), .O(new_n6548));
  inv1 g06355(.a(new_n6547), .O(new_n6549));
  nor2 g06356(.a(new_n6549), .b(new_n6517), .O(new_n6550));
  nor2 g06357(.a(new_n6550), .b(new_n6548), .O(new_n6551));
  inv1 g06358(.a(new_n6551), .O(new_n6552));
  nor2 g06359(.a(new_n6552), .b(new_n6504), .O(new_n6553));
  nor2 g06360(.a(new_n6551), .b(new_n6503), .O(new_n6554));
  nor2 g06361(.a(new_n6554), .b(new_n6553), .O(new_n6555));
  inv1 g06362(.a(new_n6555), .O(new_n6556));
  nor2 g06363(.a(new_n2433), .b(new_n1199), .O(new_n6557));
  inv1 g06364(.a(new_n6557), .O(new_n6558));
  nor2 g06365(.a(new_n2184), .b(new_n1297), .O(new_n6559));
  nor2 g06366(.a(new_n6559), .b(new_n6253), .O(new_n6560));
  nor2 g06367(.a(new_n2184), .b(new_n1425), .O(new_n6561));
  inv1 g06368(.a(new_n6561), .O(new_n6562));
  nor2 g06369(.a(new_n6562), .b(new_n6025), .O(new_n6563));
  nor2 g06370(.a(new_n6563), .b(new_n6560), .O(new_n6564));
  nor2 g06371(.a(new_n6564), .b(new_n6558), .O(new_n6565));
  inv1 g06372(.a(new_n6564), .O(new_n6566));
  nor2 g06373(.a(new_n6566), .b(new_n6557), .O(new_n6567));
  nor2 g06374(.a(new_n6567), .b(new_n6565), .O(new_n6568));
  inv1 g06375(.a(new_n6568), .O(new_n6569));
  inv1 g06376(.a(\a[47] ), .O(new_n6570));
  nor2 g06377(.a(new_n6570), .b(new_n198), .O(new_n6571));
  nor2 g06378(.a(new_n5971), .b(new_n196), .O(new_n6572));
  nor2 g06379(.a(new_n6572), .b(new_n6571), .O(new_n6573));
  nor2 g06380(.a(new_n6570), .b(new_n196), .O(new_n6574));
  inv1 g06381(.a(new_n6574), .O(new_n6575));
  nor2 g06382(.a(new_n6575), .b(new_n5982), .O(new_n6576));
  nor2 g06383(.a(new_n6576), .b(new_n6573), .O(new_n6577));
  inv1 g06384(.a(new_n6577), .O(new_n6578));
  nor2 g06385(.a(new_n6578), .b(new_n6344), .O(new_n6579));
  inv1 g06386(.a(new_n6344), .O(new_n6580));
  nor2 g06387(.a(new_n6577), .b(new_n6580), .O(new_n6581));
  nor2 g06388(.a(new_n6581), .b(new_n6579), .O(new_n6582));
  nor2 g06389(.a(new_n2826), .b(new_n847), .O(new_n6583));
  inv1 g06390(.a(new_n6583), .O(new_n6584));
  nor2 g06391(.a(new_n2660), .b(new_n941), .O(new_n6585));
  nor2 g06392(.a(new_n6585), .b(new_n6230), .O(new_n6586));
  nor2 g06393(.a(new_n2660), .b(new_n1086), .O(new_n6587));
  inv1 g06394(.a(new_n6587), .O(new_n6588));
  nor2 g06395(.a(new_n6588), .b(new_n5679), .O(new_n6589));
  nor2 g06396(.a(new_n6589), .b(new_n6586), .O(new_n6590));
  nor2 g06397(.a(new_n6590), .b(new_n6584), .O(new_n6591));
  inv1 g06398(.a(new_n6590), .O(new_n6592));
  nor2 g06399(.a(new_n6592), .b(new_n6583), .O(new_n6593));
  nor2 g06400(.a(new_n6593), .b(new_n6591), .O(new_n6594));
  nor2 g06401(.a(new_n6594), .b(new_n6582), .O(new_n6595));
  inv1 g06402(.a(new_n6582), .O(new_n6596));
  inv1 g06403(.a(new_n6594), .O(new_n6597));
  nor2 g06404(.a(new_n6597), .b(new_n6596), .O(new_n6598));
  nor2 g06405(.a(new_n6598), .b(new_n6595), .O(new_n6599));
  nor2 g06406(.a(new_n6599), .b(new_n6569), .O(new_n6600));
  inv1 g06407(.a(new_n6599), .O(new_n6601));
  nor2 g06408(.a(new_n6601), .b(new_n6568), .O(new_n6602));
  nor2 g06409(.a(new_n6602), .b(new_n6600), .O(new_n6603));
  inv1 g06410(.a(new_n6603), .O(new_n6604));
  nor2 g06411(.a(new_n6604), .b(new_n6556), .O(new_n6605));
  nor2 g06412(.a(new_n6603), .b(new_n6555), .O(new_n6606));
  nor2 g06413(.a(new_n6606), .b(new_n6605), .O(new_n6607));
  inv1 g06414(.a(new_n6607), .O(new_n6608));
  nor2 g06415(.a(new_n6244), .b(new_n6238), .O(new_n6609));
  inv1 g06416(.a(new_n6609), .O(new_n6610));
  nor2 g06417(.a(new_n6336), .b(new_n6330), .O(new_n6611));
  inv1 g06418(.a(new_n6611), .O(new_n6612));
  nor2 g06419(.a(new_n6612), .b(new_n6610), .O(new_n6613));
  nor2 g06420(.a(new_n6611), .b(new_n6609), .O(new_n6614));
  nor2 g06421(.a(new_n6614), .b(new_n6613), .O(new_n6615));
  inv1 g06422(.a(new_n6615), .O(new_n6616));
  nor2 g06423(.a(new_n6274), .b(new_n194), .O(new_n6617));
  nor2 g06424(.a(new_n6617), .b(\a[24] ), .O(new_n6618));
  nor2 g06425(.a(new_n6274), .b(new_n1736), .O(new_n6619));
  inv1 g06426(.a(new_n6619), .O(new_n6620));
  nor2 g06427(.a(new_n6620), .b(new_n194), .O(new_n6621));
  nor2 g06428(.a(new_n6621), .b(new_n6618), .O(new_n6622));
  inv1 g06429(.a(new_n6622), .O(new_n6623));
  nor2 g06430(.a(new_n6270), .b(new_n6263), .O(new_n6624));
  inv1 g06431(.a(new_n6624), .O(new_n6625));
  nor2 g06432(.a(new_n6625), .b(new_n6623), .O(new_n6626));
  nor2 g06433(.a(new_n6624), .b(new_n6622), .O(new_n6627));
  nor2 g06434(.a(new_n6627), .b(new_n6626), .O(new_n6628));
  inv1 g06435(.a(new_n6628), .O(new_n6629));
  nor2 g06436(.a(new_n6222), .b(new_n6215), .O(new_n6630));
  inv1 g06437(.a(new_n6630), .O(new_n6631));
  nor2 g06438(.a(new_n6631), .b(new_n6629), .O(new_n6632));
  nor2 g06439(.a(new_n6630), .b(new_n6628), .O(new_n6633));
  nor2 g06440(.a(new_n6633), .b(new_n6632), .O(new_n6634));
  inv1 g06441(.a(new_n6634), .O(new_n6635));
  nor2 g06442(.a(new_n6635), .b(new_n6616), .O(new_n6636));
  nor2 g06443(.a(new_n6634), .b(new_n6615), .O(new_n6637));
  nor2 g06444(.a(new_n6637), .b(new_n6636), .O(new_n6638));
  inv1 g06445(.a(new_n6638), .O(new_n6639));
  nor2 g06446(.a(new_n6639), .b(new_n6608), .O(new_n6640));
  nor2 g06447(.a(new_n6638), .b(new_n6607), .O(new_n6641));
  nor2 g06448(.a(new_n6641), .b(new_n6640), .O(new_n6642));
  inv1 g06449(.a(new_n6642), .O(new_n6643));
  nor2 g06450(.a(new_n6643), .b(new_n6479), .O(new_n6644));
  nor2 g06451(.a(new_n6642), .b(new_n6478), .O(new_n6645));
  nor2 g06452(.a(new_n6645), .b(new_n6644), .O(new_n6646));
  inv1 g06453(.a(new_n6646), .O(new_n6647));
  nor2 g06454(.a(new_n6647), .b(new_n6441), .O(new_n6648));
  inv1 g06455(.a(new_n6441), .O(new_n6649));
  nor2 g06456(.a(new_n6646), .b(new_n6649), .O(new_n6650));
  nor2 g06457(.a(new_n6650), .b(new_n6648), .O(new_n6651));
  inv1 g06458(.a(new_n6651), .O(new_n6652));
  nor2 g06459(.a(new_n6652), .b(new_n6440), .O(new_n6653));
  nor2 g06460(.a(new_n6651), .b(new_n6439), .O(new_n6654));
  nor2 g06461(.a(new_n6654), .b(new_n6653), .O(new_n6655));
  inv1 g06462(.a(new_n6655), .O(new_n6656));
  nor2 g06463(.a(new_n6656), .b(new_n6390), .O(new_n6657));
  inv1 g06464(.a(new_n6390), .O(new_n6658));
  nor2 g06465(.a(new_n6655), .b(new_n6658), .O(new_n6659));
  nor2 g06466(.a(new_n6659), .b(new_n6657), .O(new_n6660));
  inv1 g06467(.a(new_n6660), .O(new_n6661));
  nor2 g06468(.a(new_n6385), .b(new_n6378), .O(new_n6662));
  nor2 g06469(.a(new_n6662), .b(new_n6661), .O(new_n6663));
  inv1 g06470(.a(new_n6662), .O(new_n6664));
  nor2 g06471(.a(new_n6664), .b(new_n6660), .O(new_n6665));
  nor2 g06472(.a(new_n6665), .b(new_n6663), .O(new_n6666));
  inv1 g06473(.a(new_n6666), .O(\asquared[48] ));
  nor2 g06474(.a(new_n6653), .b(new_n6648), .O(new_n6668));
  inv1 g06475(.a(new_n6668), .O(new_n6669));
  nor2 g06476(.a(new_n6437), .b(new_n6396), .O(new_n6670));
  inv1 g06477(.a(new_n6670), .O(new_n6671));
  nor2 g06478(.a(new_n6433), .b(new_n6427), .O(new_n6672));
  nor2 g06479(.a(new_n6477), .b(new_n6471), .O(new_n6673));
  nor2 g06480(.a(new_n6465), .b(new_n6458), .O(new_n6674));
  inv1 g06481(.a(new_n6674), .O(new_n6675));
  nor2 g06482(.a(new_n4425), .b(new_n363), .O(new_n6676));
  inv1 g06483(.a(new_n6676), .O(new_n6677));
  nor2 g06484(.a(new_n4366), .b(new_n438), .O(new_n6678));
  nor2 g06485(.a(new_n6678), .b(new_n5665), .O(new_n6679));
  nor2 g06486(.a(new_n6531), .b(new_n6523), .O(new_n6680));
  nor2 g06487(.a(new_n6680), .b(new_n6679), .O(new_n6681));
  nor2 g06488(.a(new_n6681), .b(new_n6677), .O(new_n6682));
  inv1 g06489(.a(new_n6681), .O(new_n6683));
  nor2 g06490(.a(new_n6683), .b(new_n6676), .O(new_n6684));
  nor2 g06491(.a(new_n6684), .b(new_n6682), .O(new_n6685));
  nor2 g06492(.a(new_n3533), .b(new_n699), .O(new_n6686));
  inv1 g06493(.a(new_n6686), .O(new_n6687));
  nor2 g06494(.a(new_n5178), .b(new_n257), .O(new_n6688));
  nor2 g06495(.a(new_n3722), .b(new_n613), .O(new_n6689));
  nor2 g06496(.a(new_n6689), .b(new_n6688), .O(new_n6690));
  inv1 g06497(.a(new_n6688), .O(new_n6691));
  inv1 g06498(.a(new_n6689), .O(new_n6692));
  nor2 g06499(.a(new_n6692), .b(new_n6691), .O(new_n6693));
  nor2 g06500(.a(new_n6693), .b(new_n6690), .O(new_n6694));
  nor2 g06501(.a(new_n6694), .b(new_n6687), .O(new_n6695));
  inv1 g06502(.a(new_n6694), .O(new_n6696));
  nor2 g06503(.a(new_n6696), .b(new_n6686), .O(new_n6697));
  nor2 g06504(.a(new_n6697), .b(new_n6695), .O(new_n6698));
  nor2 g06505(.a(new_n4954), .b(new_n295), .O(new_n6699));
  inv1 g06506(.a(new_n6699), .O(new_n6700));
  nor2 g06507(.a(new_n3870), .b(new_n569), .O(new_n6701));
  nor2 g06508(.a(new_n4682), .b(new_n322), .O(new_n6702));
  nor2 g06509(.a(new_n6702), .b(new_n6701), .O(new_n6703));
  nor2 g06510(.a(new_n6451), .b(new_n5723), .O(new_n6704));
  nor2 g06511(.a(new_n6704), .b(new_n6703), .O(new_n6705));
  nor2 g06512(.a(new_n6705), .b(new_n6700), .O(new_n6706));
  inv1 g06513(.a(new_n6705), .O(new_n6707));
  nor2 g06514(.a(new_n6707), .b(new_n6699), .O(new_n6708));
  nor2 g06515(.a(new_n6708), .b(new_n6706), .O(new_n6709));
  nor2 g06516(.a(new_n6709), .b(new_n6698), .O(new_n6710));
  inv1 g06517(.a(new_n6698), .O(new_n6711));
  inv1 g06518(.a(new_n6709), .O(new_n6712));
  nor2 g06519(.a(new_n6712), .b(new_n6711), .O(new_n6713));
  nor2 g06520(.a(new_n6713), .b(new_n6710), .O(new_n6714));
  inv1 g06521(.a(new_n6714), .O(new_n6715));
  nor2 g06522(.a(new_n6715), .b(new_n6685), .O(new_n6716));
  inv1 g06523(.a(new_n6685), .O(new_n6717));
  nor2 g06524(.a(new_n6714), .b(new_n6717), .O(new_n6718));
  nor2 g06525(.a(new_n6718), .b(new_n6716), .O(new_n6719));
  nor2 g06526(.a(new_n6719), .b(new_n6675), .O(new_n6720));
  inv1 g06527(.a(new_n6719), .O(new_n6721));
  nor2 g06528(.a(new_n6721), .b(new_n6674), .O(new_n6722));
  nor2 g06529(.a(new_n6722), .b(new_n6720), .O(new_n6723));
  nor2 g06530(.a(new_n2826), .b(new_n941), .O(new_n6724));
  inv1 g06531(.a(new_n6724), .O(new_n6725));
  nor2 g06532(.a(new_n2506), .b(new_n1199), .O(new_n6726));
  nor2 g06533(.a(new_n6726), .b(new_n6587), .O(new_n6727));
  nor2 g06534(.a(new_n2660), .b(new_n1199), .O(new_n6728));
  inv1 g06535(.a(new_n6728), .O(new_n6729));
  nor2 g06536(.a(new_n6729), .b(new_n6231), .O(new_n6730));
  nor2 g06537(.a(new_n6730), .b(new_n6727), .O(new_n6731));
  nor2 g06538(.a(new_n6731), .b(new_n6725), .O(new_n6732));
  inv1 g06539(.a(new_n6731), .O(new_n6733));
  nor2 g06540(.a(new_n6733), .b(new_n6724), .O(new_n6734));
  nor2 g06541(.a(new_n6734), .b(new_n6732), .O(new_n6735));
  inv1 g06542(.a(new_n6735), .O(new_n6736));
  nor2 g06543(.a(new_n5796), .b(new_n214), .O(new_n6737));
  nor2 g06544(.a(new_n5393), .b(new_n229), .O(new_n6738));
  nor2 g06545(.a(new_n3231), .b(new_n800), .O(new_n6739));
  nor2 g06546(.a(new_n6739), .b(new_n6738), .O(new_n6740));
  nor2 g06547(.a(new_n6493), .b(new_n4248), .O(new_n6741));
  nor2 g06548(.a(new_n6741), .b(new_n6740), .O(new_n6742));
  inv1 g06549(.a(new_n6742), .O(new_n6743));
  nor2 g06550(.a(new_n6743), .b(new_n6737), .O(new_n6744));
  inv1 g06551(.a(new_n6737), .O(new_n6745));
  nor2 g06552(.a(new_n6742), .b(new_n6745), .O(new_n6746));
  nor2 g06553(.a(new_n6746), .b(new_n6744), .O(new_n6747));
  nor2 g06554(.a(new_n2433), .b(new_n1297), .O(new_n6748));
  inv1 g06555(.a(new_n6748), .O(new_n6749));
  nor2 g06556(.a(new_n2121), .b(new_n1493), .O(new_n6750));
  nor2 g06557(.a(new_n6750), .b(new_n6561), .O(new_n6751));
  nor2 g06558(.a(new_n2184), .b(new_n1493), .O(new_n6752));
  inv1 g06559(.a(new_n6752), .O(new_n6753));
  nor2 g06560(.a(new_n6753), .b(new_n6254), .O(new_n6754));
  nor2 g06561(.a(new_n6754), .b(new_n6751), .O(new_n6755));
  nor2 g06562(.a(new_n6755), .b(new_n6749), .O(new_n6756));
  inv1 g06563(.a(new_n6755), .O(new_n6757));
  nor2 g06564(.a(new_n6757), .b(new_n6748), .O(new_n6758));
  nor2 g06565(.a(new_n6758), .b(new_n6756), .O(new_n6759));
  nor2 g06566(.a(new_n6759), .b(new_n6747), .O(new_n6760));
  inv1 g06567(.a(new_n6747), .O(new_n6761));
  inv1 g06568(.a(new_n6759), .O(new_n6762));
  nor2 g06569(.a(new_n6762), .b(new_n6761), .O(new_n6763));
  nor2 g06570(.a(new_n6763), .b(new_n6760), .O(new_n6764));
  nor2 g06571(.a(new_n6764), .b(new_n6736), .O(new_n6765));
  inv1 g06572(.a(new_n6764), .O(new_n6766));
  nor2 g06573(.a(new_n6766), .b(new_n6735), .O(new_n6767));
  nor2 g06574(.a(new_n6767), .b(new_n6765), .O(new_n6768));
  nor2 g06575(.a(new_n6768), .b(new_n6723), .O(new_n6769));
  inv1 g06576(.a(new_n6723), .O(new_n6770));
  inv1 g06577(.a(new_n6768), .O(new_n6771));
  nor2 g06578(.a(new_n6771), .b(new_n6770), .O(new_n6772));
  nor2 g06579(.a(new_n6772), .b(new_n6769), .O(new_n6773));
  inv1 g06580(.a(new_n6773), .O(new_n6774));
  nor2 g06581(.a(new_n6774), .b(new_n6673), .O(new_n6775));
  inv1 g06582(.a(new_n6673), .O(new_n6776));
  nor2 g06583(.a(new_n6773), .b(new_n6776), .O(new_n6777));
  nor2 g06584(.a(new_n6777), .b(new_n6775), .O(new_n6778));
  inv1 g06585(.a(new_n6778), .O(new_n6779));
  nor2 g06586(.a(new_n6779), .b(new_n6672), .O(new_n6780));
  inv1 g06587(.a(new_n6672), .O(new_n6781));
  nor2 g06588(.a(new_n6778), .b(new_n6781), .O(new_n6782));
  nor2 g06589(.a(new_n6782), .b(new_n6780), .O(new_n6783));
  nor2 g06590(.a(new_n6783), .b(new_n6671), .O(new_n6784));
  inv1 g06591(.a(new_n6783), .O(new_n6785));
  nor2 g06592(.a(new_n6785), .b(new_n6670), .O(new_n6786));
  nor2 g06593(.a(new_n6786), .b(new_n6784), .O(new_n6787));
  inv1 g06594(.a(new_n6787), .O(new_n6788));
  nor2 g06595(.a(new_n6567), .b(new_n6560), .O(new_n6789));
  nor2 g06596(.a(new_n6527), .b(new_n6520), .O(new_n6790));
  nor2 g06597(.a(new_n6790), .b(new_n6789), .O(new_n6791));
  inv1 g06598(.a(new_n6789), .O(new_n6792));
  inv1 g06599(.a(new_n6790), .O(new_n6793));
  nor2 g06600(.a(new_n6793), .b(new_n6792), .O(new_n6794));
  nor2 g06601(.a(new_n6794), .b(new_n6791), .O(new_n6795));
  nor2 g06602(.a(new_n6516), .b(new_n6509), .O(new_n6796));
  nor2 g06603(.a(new_n6796), .b(new_n6795), .O(new_n6797));
  inv1 g06604(.a(new_n6795), .O(new_n6798));
  inv1 g06605(.a(new_n6796), .O(new_n6799));
  nor2 g06606(.a(new_n6799), .b(new_n6798), .O(new_n6800));
  nor2 g06607(.a(new_n6800), .b(new_n6797), .O(new_n6801));
  nor2 g06608(.a(new_n6550), .b(new_n6543), .O(new_n6802));
  inv1 g06609(.a(new_n6802), .O(new_n6803));
  nor2 g06610(.a(new_n6803), .b(new_n6801), .O(new_n6804));
  inv1 g06611(.a(new_n6801), .O(new_n6805));
  nor2 g06612(.a(new_n6802), .b(new_n6805), .O(new_n6806));
  nor2 g06613(.a(new_n6806), .b(new_n6804), .O(new_n6807));
  nor2 g06614(.a(new_n6456), .b(new_n6449), .O(new_n6808));
  nor2 g06615(.a(new_n6541), .b(new_n6534), .O(new_n6809));
  nor2 g06616(.a(new_n6809), .b(new_n6808), .O(new_n6810));
  inv1 g06617(.a(new_n6808), .O(new_n6811));
  inv1 g06618(.a(new_n6809), .O(new_n6812));
  nor2 g06619(.a(new_n6812), .b(new_n6811), .O(new_n6813));
  nor2 g06620(.a(new_n6813), .b(new_n6810), .O(new_n6814));
  inv1 g06621(.a(new_n6814), .O(new_n6815));
  nor2 g06622(.a(new_n6274), .b(new_n196), .O(new_n6816));
  inv1 g06623(.a(new_n6816), .O(new_n6817));
  nor2 g06624(.a(new_n5971), .b(new_n203), .O(new_n6818));
  nor2 g06625(.a(new_n3057), .b(new_n847), .O(new_n6819));
  nor2 g06626(.a(new_n6819), .b(new_n6818), .O(new_n6820));
  inv1 g06627(.a(new_n6818), .O(new_n6821));
  inv1 g06628(.a(new_n6819), .O(new_n6822));
  nor2 g06629(.a(new_n6822), .b(new_n6821), .O(new_n6823));
  nor2 g06630(.a(new_n6823), .b(new_n6820), .O(new_n6824));
  nor2 g06631(.a(new_n6824), .b(new_n6817), .O(new_n6825));
  inv1 g06632(.a(new_n6824), .O(new_n6826));
  nor2 g06633(.a(new_n6826), .b(new_n6816), .O(new_n6827));
  nor2 g06634(.a(new_n6827), .b(new_n6825), .O(new_n6828));
  nor2 g06635(.a(new_n6828), .b(new_n6815), .O(new_n6829));
  inv1 g06636(.a(new_n6828), .O(new_n6830));
  nor2 g06637(.a(new_n6830), .b(new_n6814), .O(new_n6831));
  nor2 g06638(.a(new_n6831), .b(new_n6829), .O(new_n6832));
  nor2 g06639(.a(new_n6832), .b(new_n6807), .O(new_n6833));
  inv1 g06640(.a(new_n6807), .O(new_n6834));
  inv1 g06641(.a(new_n6832), .O(new_n6835));
  nor2 g06642(.a(new_n6835), .b(new_n6834), .O(new_n6836));
  nor2 g06643(.a(new_n6836), .b(new_n6833), .O(new_n6837));
  inv1 g06644(.a(new_n6837), .O(new_n6838));
  nor2 g06645(.a(new_n6605), .b(new_n6553), .O(new_n6839));
  nor2 g06646(.a(new_n6839), .b(new_n6838), .O(new_n6840));
  inv1 g06647(.a(new_n6839), .O(new_n6841));
  nor2 g06648(.a(new_n6841), .b(new_n6837), .O(new_n6842));
  nor2 g06649(.a(new_n6842), .b(new_n6840), .O(new_n6843));
  inv1 g06650(.a(new_n6843), .O(new_n6844));
  nor2 g06651(.a(new_n6593), .b(new_n6586), .O(new_n6845));
  nor2 g06652(.a(new_n6498), .b(new_n6491), .O(new_n6846));
  nor2 g06653(.a(new_n6846), .b(new_n6845), .O(new_n6847));
  inv1 g06654(.a(new_n6845), .O(new_n6848));
  inv1 g06655(.a(new_n6846), .O(new_n6849));
  nor2 g06656(.a(new_n6849), .b(new_n6848), .O(new_n6850));
  nor2 g06657(.a(new_n6850), .b(new_n6847), .O(new_n6851));
  nor2 g06658(.a(new_n6579), .b(new_n6573), .O(new_n6852));
  nor2 g06659(.a(new_n6852), .b(new_n6851), .O(new_n6853));
  inv1 g06660(.a(new_n6851), .O(new_n6854));
  inv1 g06661(.a(new_n6852), .O(new_n6855));
  nor2 g06662(.a(new_n6855), .b(new_n6854), .O(new_n6856));
  nor2 g06663(.a(new_n6856), .b(new_n6853), .O(new_n6857));
  inv1 g06664(.a(new_n6857), .O(new_n6858));
  nor2 g06665(.a(new_n6632), .b(new_n6626), .O(new_n6859));
  inv1 g06666(.a(new_n6859), .O(new_n6860));
  nor2 g06667(.a(new_n6602), .b(new_n6595), .O(new_n6861));
  inv1 g06668(.a(new_n6861), .O(new_n6862));
  nor2 g06669(.a(new_n6862), .b(new_n6860), .O(new_n6863));
  nor2 g06670(.a(new_n6861), .b(new_n6859), .O(new_n6864));
  nor2 g06671(.a(new_n6864), .b(new_n6863), .O(new_n6865));
  inv1 g06672(.a(new_n6865), .O(new_n6866));
  nor2 g06673(.a(new_n6866), .b(new_n6858), .O(new_n6867));
  nor2 g06674(.a(new_n6865), .b(new_n6857), .O(new_n6868));
  nor2 g06675(.a(new_n6868), .b(new_n6867), .O(new_n6869));
  inv1 g06676(.a(new_n6869), .O(new_n6870));
  nor2 g06677(.a(new_n6870), .b(new_n6844), .O(new_n6871));
  nor2 g06678(.a(new_n6869), .b(new_n6843), .O(new_n6872));
  nor2 g06679(.a(new_n6872), .b(new_n6871), .O(new_n6873));
  inv1 g06680(.a(new_n6873), .O(new_n6874));
  nor2 g06681(.a(new_n6644), .b(new_n6640), .O(new_n6875));
  nor2 g06682(.a(new_n6422), .b(new_n6416), .O(new_n6876));
  inv1 g06683(.a(new_n6876), .O(new_n6877));
  nor2 g06684(.a(new_n6636), .b(new_n6614), .O(new_n6878));
  inv1 g06685(.a(new_n6878), .O(new_n6879));
  nor2 g06686(.a(new_n6879), .b(new_n6877), .O(new_n6880));
  nor2 g06687(.a(new_n6878), .b(new_n6876), .O(new_n6881));
  nor2 g06688(.a(new_n6881), .b(new_n6880), .O(new_n6882));
  inv1 g06689(.a(new_n6882), .O(new_n6883));
  nor2 g06690(.a(new_n6410), .b(new_n6404), .O(new_n6884));
  inv1 g06691(.a(new_n6884), .O(new_n6885));
  nor2 g06692(.a(new_n6570), .b(new_n194), .O(new_n6886));
  nor2 g06693(.a(new_n6886), .b(new_n6535), .O(new_n6887));
  inv1 g06694(.a(new_n6886), .O(new_n6888));
  nor2 g06695(.a(new_n6888), .b(new_n6536), .O(new_n6889));
  nor2 g06696(.a(new_n6889), .b(new_n6887), .O(new_n6890));
  inv1 g06697(.a(new_n6890), .O(new_n6891));
  inv1 g06698(.a(new_n6621), .O(new_n6892));
  inv1 g06699(.a(\a[48] ), .O(new_n6893));
  nor2 g06700(.a(new_n6893), .b(new_n198), .O(new_n6894));
  inv1 g06701(.a(new_n6894), .O(new_n6895));
  nor2 g06702(.a(new_n6895), .b(new_n6892), .O(new_n6896));
  nor2 g06703(.a(new_n6894), .b(new_n6621), .O(new_n6897));
  nor2 g06704(.a(new_n6897), .b(new_n6896), .O(new_n6898));
  inv1 g06705(.a(new_n6898), .O(new_n6899));
  nor2 g06706(.a(new_n6899), .b(new_n6891), .O(new_n6900));
  nor2 g06707(.a(new_n6898), .b(new_n6890), .O(new_n6901));
  nor2 g06708(.a(new_n6901), .b(new_n6900), .O(new_n6902));
  nor2 g06709(.a(new_n6902), .b(new_n6885), .O(new_n6903));
  inv1 g06710(.a(new_n6902), .O(new_n6904));
  nor2 g06711(.a(new_n6904), .b(new_n6884), .O(new_n6905));
  nor2 g06712(.a(new_n6905), .b(new_n6903), .O(new_n6906));
  nor2 g06713(.a(new_n6500), .b(new_n6485), .O(new_n6907));
  inv1 g06714(.a(new_n6907), .O(new_n6908));
  nor2 g06715(.a(new_n6908), .b(new_n6906), .O(new_n6909));
  inv1 g06716(.a(new_n6906), .O(new_n6910));
  nor2 g06717(.a(new_n6907), .b(new_n6910), .O(new_n6911));
  nor2 g06718(.a(new_n6911), .b(new_n6909), .O(new_n6912));
  inv1 g06719(.a(new_n6912), .O(new_n6913));
  nor2 g06720(.a(new_n6913), .b(new_n6883), .O(new_n6914));
  nor2 g06721(.a(new_n6912), .b(new_n6882), .O(new_n6915));
  nor2 g06722(.a(new_n6915), .b(new_n6914), .O(new_n6916));
  inv1 g06723(.a(new_n6916), .O(new_n6917));
  nor2 g06724(.a(new_n6917), .b(new_n6875), .O(new_n6918));
  inv1 g06725(.a(new_n6875), .O(new_n6919));
  nor2 g06726(.a(new_n6916), .b(new_n6919), .O(new_n6920));
  nor2 g06727(.a(new_n6920), .b(new_n6918), .O(new_n6921));
  inv1 g06728(.a(new_n6921), .O(new_n6922));
  nor2 g06729(.a(new_n6922), .b(new_n6874), .O(new_n6923));
  nor2 g06730(.a(new_n6921), .b(new_n6873), .O(new_n6924));
  nor2 g06731(.a(new_n6924), .b(new_n6923), .O(new_n6925));
  inv1 g06732(.a(new_n6925), .O(new_n6926));
  nor2 g06733(.a(new_n6926), .b(new_n6788), .O(new_n6927));
  nor2 g06734(.a(new_n6925), .b(new_n6787), .O(new_n6928));
  nor2 g06735(.a(new_n6928), .b(new_n6927), .O(new_n6929));
  nor2 g06736(.a(new_n6929), .b(new_n6669), .O(new_n6930));
  inv1 g06737(.a(new_n6929), .O(new_n6931));
  nor2 g06738(.a(new_n6931), .b(new_n6668), .O(new_n6932));
  nor2 g06739(.a(new_n6932), .b(new_n6930), .O(new_n6933));
  inv1 g06740(.a(new_n6933), .O(new_n6934));
  nor2 g06741(.a(new_n6663), .b(new_n6659), .O(new_n6935));
  nor2 g06742(.a(new_n6935), .b(new_n6934), .O(new_n6936));
  inv1 g06743(.a(new_n6935), .O(new_n6937));
  nor2 g06744(.a(new_n6937), .b(new_n6933), .O(new_n6938));
  nor2 g06745(.a(new_n6938), .b(new_n6936), .O(new_n6939));
  inv1 g06746(.a(new_n6939), .O(\asquared[49] ));
  nor2 g06747(.a(new_n6923), .b(new_n6918), .O(new_n6941));
  nor2 g06748(.a(new_n6871), .b(new_n6840), .O(new_n6942));
  nor2 g06749(.a(new_n6914), .b(new_n6881), .O(new_n6943));
  nor2 g06750(.a(new_n3231), .b(new_n847), .O(new_n6944));
  inv1 g06751(.a(new_n6944), .O(new_n6945));
  nor2 g06752(.a(new_n3057), .b(new_n941), .O(new_n6946));
  nor2 g06753(.a(new_n2826), .b(new_n1086), .O(new_n6947));
  nor2 g06754(.a(new_n6947), .b(new_n6946), .O(new_n6948));
  nor2 g06755(.a(new_n3057), .b(new_n1086), .O(new_n6949));
  inv1 g06756(.a(new_n6949), .O(new_n6950));
  nor2 g06757(.a(new_n6950), .b(new_n6725), .O(new_n6951));
  nor2 g06758(.a(new_n6951), .b(new_n6948), .O(new_n6952));
  nor2 g06759(.a(new_n6952), .b(new_n6945), .O(new_n6953));
  inv1 g06760(.a(new_n6952), .O(new_n6954));
  nor2 g06761(.a(new_n6954), .b(new_n6944), .O(new_n6955));
  nor2 g06762(.a(new_n6955), .b(new_n6953), .O(new_n6956));
  nor2 g06763(.a(new_n6900), .b(new_n6896), .O(new_n6957));
  inv1 g06764(.a(\a[49] ), .O(new_n6958));
  nor2 g06765(.a(new_n6958), .b(new_n198), .O(new_n6959));
  inv1 g06766(.a(new_n6959), .O(new_n6960));
  nor2 g06767(.a(new_n5971), .b(new_n214), .O(new_n6961));
  nor2 g06768(.a(new_n5796), .b(new_n229), .O(new_n6962));
  nor2 g06769(.a(new_n6962), .b(new_n6961), .O(new_n6963));
  nor2 g06770(.a(new_n5971), .b(new_n229), .O(new_n6964));
  inv1 g06771(.a(new_n6964), .O(new_n6965));
  nor2 g06772(.a(new_n6965), .b(new_n6745), .O(new_n6966));
  nor2 g06773(.a(new_n6966), .b(new_n6963), .O(new_n6967));
  nor2 g06774(.a(new_n6967), .b(new_n6960), .O(new_n6968));
  inv1 g06775(.a(new_n6967), .O(new_n6969));
  nor2 g06776(.a(new_n6969), .b(new_n6959), .O(new_n6970));
  nor2 g06777(.a(new_n6970), .b(new_n6968), .O(new_n6971));
  nor2 g06778(.a(new_n6971), .b(new_n6957), .O(new_n6972));
  inv1 g06779(.a(new_n6957), .O(new_n6973));
  inv1 g06780(.a(new_n6971), .O(new_n6974));
  nor2 g06781(.a(new_n6974), .b(new_n6973), .O(new_n6975));
  nor2 g06782(.a(new_n6975), .b(new_n6972), .O(new_n6976));
  inv1 g06783(.a(new_n6976), .O(new_n6977));
  nor2 g06784(.a(new_n6977), .b(new_n6956), .O(new_n6978));
  inv1 g06785(.a(new_n6956), .O(new_n6979));
  nor2 g06786(.a(new_n6976), .b(new_n6979), .O(new_n6980));
  nor2 g06787(.a(new_n6980), .b(new_n6978), .O(new_n6981));
  inv1 g06788(.a(new_n6981), .O(new_n6982));
  nor2 g06789(.a(new_n4682), .b(new_n363), .O(new_n6983));
  inv1 g06790(.a(new_n6983), .O(new_n6984));
  nor2 g06791(.a(new_n4093), .b(new_n569), .O(new_n6985));
  nor2 g06792(.a(new_n4425), .b(new_n438), .O(new_n6986));
  nor2 g06793(.a(new_n6986), .b(new_n6985), .O(new_n6987));
  nor2 g06794(.a(new_n4425), .b(new_n569), .O(new_n6988));
  inv1 g06795(.a(new_n6988), .O(new_n6989));
  nor2 g06796(.a(new_n6989), .b(new_n6531), .O(new_n6990));
  nor2 g06797(.a(new_n6990), .b(new_n6987), .O(new_n6991));
  nor2 g06798(.a(new_n6991), .b(new_n6984), .O(new_n6992));
  inv1 g06799(.a(new_n6991), .O(new_n6993));
  nor2 g06800(.a(new_n6993), .b(new_n6983), .O(new_n6994));
  nor2 g06801(.a(new_n6994), .b(new_n6992), .O(new_n6995));
  inv1 g06802(.a(new_n6995), .O(new_n6996));
  nor2 g06803(.a(new_n6274), .b(new_n203), .O(new_n6997));
  nor2 g06804(.a(new_n6997), .b(new_n6574), .O(new_n6998));
  nor2 g06805(.a(new_n6570), .b(new_n203), .O(new_n6999));
  inv1 g06806(.a(new_n6999), .O(new_n7000));
  nor2 g06807(.a(new_n7000), .b(new_n6817), .O(new_n7001));
  nor2 g06808(.a(new_n7001), .b(new_n6998), .O(new_n7002));
  inv1 g06809(.a(new_n7002), .O(new_n7003));
  nor2 g06810(.a(new_n7003), .b(new_n6752), .O(new_n7004));
  nor2 g06811(.a(new_n7002), .b(new_n6753), .O(new_n7005));
  nor2 g06812(.a(new_n7005), .b(new_n7004), .O(new_n7006));
  nor2 g06813(.a(new_n2506), .b(new_n1297), .O(new_n7007));
  nor2 g06814(.a(new_n2433), .b(new_n1425), .O(new_n7008));
  nor2 g06815(.a(new_n7008), .b(new_n7007), .O(new_n7009));
  nor2 g06816(.a(new_n2506), .b(new_n1425), .O(new_n7010));
  inv1 g06817(.a(new_n7010), .O(new_n7011));
  nor2 g06818(.a(new_n7011), .b(new_n6749), .O(new_n7012));
  nor2 g06819(.a(new_n7012), .b(new_n7009), .O(new_n7013));
  nor2 g06820(.a(new_n7013), .b(new_n6729), .O(new_n7014));
  inv1 g06821(.a(new_n7013), .O(new_n7015));
  nor2 g06822(.a(new_n7015), .b(new_n6728), .O(new_n7016));
  nor2 g06823(.a(new_n7016), .b(new_n7014), .O(new_n7017));
  nor2 g06824(.a(new_n7017), .b(new_n7006), .O(new_n7018));
  inv1 g06825(.a(new_n7006), .O(new_n7019));
  inv1 g06826(.a(new_n7017), .O(new_n7020));
  nor2 g06827(.a(new_n7020), .b(new_n7019), .O(new_n7021));
  nor2 g06828(.a(new_n7021), .b(new_n7018), .O(new_n7022));
  nor2 g06829(.a(new_n7022), .b(new_n6996), .O(new_n7023));
  inv1 g06830(.a(new_n7022), .O(new_n7024));
  nor2 g06831(.a(new_n7024), .b(new_n6995), .O(new_n7025));
  nor2 g06832(.a(new_n7025), .b(new_n7023), .O(new_n7026));
  inv1 g06833(.a(new_n7026), .O(new_n7027));
  nor2 g06834(.a(new_n7027), .b(new_n6982), .O(new_n7028));
  nor2 g06835(.a(new_n7026), .b(new_n6981), .O(new_n7029));
  nor2 g06836(.a(new_n7029), .b(new_n7028), .O(new_n7030));
  inv1 g06837(.a(new_n7030), .O(new_n7031));
  nor2 g06838(.a(new_n3533), .b(new_n800), .O(new_n7032));
  inv1 g06839(.a(new_n7032), .O(new_n7033));
  nor2 g06840(.a(new_n5393), .b(new_n257), .O(new_n7034));
  nor2 g06841(.a(new_n3722), .b(new_n699), .O(new_n7035));
  nor2 g06842(.a(new_n7035), .b(new_n7034), .O(new_n7036));
  inv1 g06843(.a(new_n5005), .O(new_n7037));
  nor2 g06844(.a(new_n5393), .b(new_n699), .O(new_n7038));
  inv1 g06845(.a(new_n7038), .O(new_n7039));
  nor2 g06846(.a(new_n7039), .b(new_n7037), .O(new_n7040));
  nor2 g06847(.a(new_n7040), .b(new_n7036), .O(new_n7041));
  nor2 g06848(.a(new_n7041), .b(new_n7033), .O(new_n7042));
  inv1 g06849(.a(new_n7041), .O(new_n7043));
  nor2 g06850(.a(new_n7043), .b(new_n7032), .O(new_n7044));
  nor2 g06851(.a(new_n7044), .b(new_n7042), .O(new_n7045));
  inv1 g06852(.a(new_n7045), .O(new_n7046));
  nor2 g06853(.a(new_n3870), .b(new_n613), .O(new_n7047));
  nor2 g06854(.a(new_n4954), .b(new_n322), .O(new_n7048));
  nor2 g06855(.a(new_n5178), .b(new_n295), .O(new_n7049));
  nor2 g06856(.a(new_n7049), .b(new_n7048), .O(new_n7050));
  nor2 g06857(.a(new_n5178), .b(new_n322), .O(new_n7051));
  inv1 g06858(.a(new_n7051), .O(new_n7052));
  nor2 g06859(.a(new_n7052), .b(new_n6700), .O(new_n7053));
  nor2 g06860(.a(new_n7053), .b(new_n7050), .O(new_n7054));
  inv1 g06861(.a(new_n7054), .O(new_n7055));
  nor2 g06862(.a(new_n7055), .b(new_n7047), .O(new_n7056));
  inv1 g06863(.a(new_n7047), .O(new_n7057));
  nor2 g06864(.a(new_n7054), .b(new_n7057), .O(new_n7058));
  nor2 g06865(.a(new_n7058), .b(new_n7056), .O(new_n7059));
  nor2 g06866(.a(new_n1903), .b(new_n1736), .O(new_n7060));
  nor2 g06867(.a(new_n2121), .b(new_n1647), .O(new_n7061));
  nor2 g06868(.a(new_n7061), .b(new_n7060), .O(new_n7062));
  inv1 g06869(.a(new_n7060), .O(new_n7063));
  inv1 g06870(.a(new_n7061), .O(new_n7064));
  nor2 g06871(.a(new_n7064), .b(new_n7063), .O(new_n7065));
  nor2 g06872(.a(new_n7065), .b(new_n7062), .O(new_n7066));
  nor2 g06873(.a(new_n7066), .b(new_n6523), .O(new_n7067));
  inv1 g06874(.a(new_n7066), .O(new_n7068));
  nor2 g06875(.a(new_n7068), .b(new_n6522), .O(new_n7069));
  nor2 g06876(.a(new_n7069), .b(new_n7067), .O(new_n7070));
  nor2 g06877(.a(new_n7070), .b(new_n7059), .O(new_n7071));
  inv1 g06878(.a(new_n7059), .O(new_n7072));
  inv1 g06879(.a(new_n7070), .O(new_n7073));
  nor2 g06880(.a(new_n7073), .b(new_n7072), .O(new_n7074));
  nor2 g06881(.a(new_n7074), .b(new_n7071), .O(new_n7075));
  nor2 g06882(.a(new_n7075), .b(new_n7046), .O(new_n7076));
  inv1 g06883(.a(new_n7075), .O(new_n7077));
  nor2 g06884(.a(new_n7077), .b(new_n7045), .O(new_n7078));
  nor2 g06885(.a(new_n7078), .b(new_n7076), .O(new_n7079));
  inv1 g06886(.a(new_n7079), .O(new_n7080));
  nor2 g06887(.a(new_n7080), .b(new_n7031), .O(new_n7081));
  nor2 g06888(.a(new_n7079), .b(new_n7030), .O(new_n7082));
  nor2 g06889(.a(new_n7082), .b(new_n7081), .O(new_n7083));
  inv1 g06890(.a(new_n7083), .O(new_n7084));
  nor2 g06891(.a(new_n7084), .b(new_n6943), .O(new_n7085));
  inv1 g06892(.a(new_n6943), .O(new_n7086));
  nor2 g06893(.a(new_n7083), .b(new_n7086), .O(new_n7087));
  nor2 g06894(.a(new_n7087), .b(new_n7085), .O(new_n7088));
  inv1 g06895(.a(new_n7088), .O(new_n7089));
  nor2 g06896(.a(new_n7089), .b(new_n6942), .O(new_n7090));
  inv1 g06897(.a(new_n6942), .O(new_n7091));
  nor2 g06898(.a(new_n7088), .b(new_n7091), .O(new_n7092));
  nor2 g06899(.a(new_n7092), .b(new_n7090), .O(new_n7093));
  inv1 g06900(.a(new_n7093), .O(new_n7094));
  nor2 g06901(.a(new_n7094), .b(new_n6941), .O(new_n7095));
  inv1 g06902(.a(new_n6941), .O(new_n7096));
  nor2 g06903(.a(new_n7093), .b(new_n7096), .O(new_n7097));
  nor2 g06904(.a(new_n7097), .b(new_n7095), .O(new_n7098));
  inv1 g06905(.a(new_n7098), .O(new_n7099));
  nor2 g06906(.a(new_n6697), .b(new_n6690), .O(new_n7100));
  nor2 g06907(.a(new_n6734), .b(new_n6727), .O(new_n7101));
  nor2 g06908(.a(new_n7101), .b(new_n7100), .O(new_n7102));
  inv1 g06909(.a(new_n7100), .O(new_n7103));
  inv1 g06910(.a(new_n7101), .O(new_n7104));
  nor2 g06911(.a(new_n7104), .b(new_n7103), .O(new_n7105));
  nor2 g06912(.a(new_n7105), .b(new_n7102), .O(new_n7106));
  nor2 g06913(.a(new_n6708), .b(new_n6703), .O(new_n7107));
  nor2 g06914(.a(new_n7107), .b(new_n7106), .O(new_n7108));
  inv1 g06915(.a(new_n7106), .O(new_n7109));
  inv1 g06916(.a(new_n7107), .O(new_n7110));
  nor2 g06917(.a(new_n7110), .b(new_n7109), .O(new_n7111));
  nor2 g06918(.a(new_n7111), .b(new_n7108), .O(new_n7112));
  nor2 g06919(.a(new_n6767), .b(new_n6760), .O(new_n7113));
  inv1 g06920(.a(new_n7113), .O(new_n7114));
  nor2 g06921(.a(new_n7114), .b(new_n7112), .O(new_n7115));
  inv1 g06922(.a(new_n7112), .O(new_n7116));
  nor2 g06923(.a(new_n7113), .b(new_n7116), .O(new_n7117));
  nor2 g06924(.a(new_n7117), .b(new_n7115), .O(new_n7118));
  nor2 g06925(.a(new_n6911), .b(new_n6905), .O(new_n7119));
  inv1 g06926(.a(new_n7119), .O(new_n7120));
  nor2 g06927(.a(new_n7120), .b(new_n7118), .O(new_n7121));
  inv1 g06928(.a(new_n7118), .O(new_n7122));
  nor2 g06929(.a(new_n7119), .b(new_n7122), .O(new_n7123));
  nor2 g06930(.a(new_n7123), .b(new_n7121), .O(new_n7124));
  inv1 g06931(.a(new_n7124), .O(new_n7125));
  nor2 g06932(.a(new_n6772), .b(new_n6722), .O(new_n7126));
  nor2 g06933(.a(new_n7126), .b(new_n7125), .O(new_n7127));
  inv1 g06934(.a(new_n7126), .O(new_n7128));
  nor2 g06935(.a(new_n7128), .b(new_n7124), .O(new_n7129));
  nor2 g06936(.a(new_n7129), .b(new_n7127), .O(new_n7130));
  inv1 g06937(.a(new_n7130), .O(new_n7131));
  nor2 g06938(.a(new_n6827), .b(new_n6820), .O(new_n7132));
  nor2 g06939(.a(new_n6744), .b(new_n6740), .O(new_n7133));
  nor2 g06940(.a(new_n7133), .b(new_n7132), .O(new_n7134));
  inv1 g06941(.a(new_n7132), .O(new_n7135));
  inv1 g06942(.a(new_n7133), .O(new_n7136));
  nor2 g06943(.a(new_n7136), .b(new_n7135), .O(new_n7137));
  nor2 g06944(.a(new_n7137), .b(new_n7134), .O(new_n7138));
  nor2 g06945(.a(new_n6758), .b(new_n6751), .O(new_n7139));
  nor2 g06946(.a(new_n7139), .b(new_n7138), .O(new_n7140));
  inv1 g06947(.a(new_n7138), .O(new_n7141));
  inv1 g06948(.a(new_n7139), .O(new_n7142));
  nor2 g06949(.a(new_n7142), .b(new_n7141), .O(new_n7143));
  nor2 g06950(.a(new_n7143), .b(new_n7140), .O(new_n7144));
  inv1 g06951(.a(new_n7144), .O(new_n7145));
  nor2 g06952(.a(new_n6716), .b(new_n6710), .O(new_n7146));
  nor2 g06953(.a(new_n2017), .b(new_n6893), .O(new_n7147));
  nor2 g06954(.a(new_n6893), .b(new_n194), .O(new_n7148));
  nor2 g06955(.a(new_n7148), .b(\a[25] ), .O(new_n7149));
  nor2 g06956(.a(new_n7149), .b(new_n7147), .O(new_n7150));
  nor2 g06957(.a(new_n7150), .b(new_n6889), .O(new_n7151));
  inv1 g06958(.a(new_n6889), .O(new_n7152));
  nor2 g06959(.a(new_n7152), .b(\a[48] ), .O(new_n7153));
  nor2 g06960(.a(new_n7153), .b(new_n7151), .O(new_n7154));
  inv1 g06961(.a(new_n7154), .O(new_n7155));
  nor2 g06962(.a(new_n6684), .b(new_n6679), .O(new_n7156));
  inv1 g06963(.a(new_n7156), .O(new_n7157));
  nor2 g06964(.a(new_n7157), .b(new_n7155), .O(new_n7158));
  nor2 g06965(.a(new_n7156), .b(new_n7154), .O(new_n7159));
  nor2 g06966(.a(new_n7159), .b(new_n7158), .O(new_n7160));
  inv1 g06967(.a(new_n7160), .O(new_n7161));
  nor2 g06968(.a(new_n7161), .b(new_n7146), .O(new_n7162));
  inv1 g06969(.a(new_n7146), .O(new_n7163));
  nor2 g06970(.a(new_n7160), .b(new_n7163), .O(new_n7164));
  nor2 g06971(.a(new_n7164), .b(new_n7162), .O(new_n7165));
  inv1 g06972(.a(new_n7165), .O(new_n7166));
  nor2 g06973(.a(new_n7166), .b(new_n7145), .O(new_n7167));
  nor2 g06974(.a(new_n7165), .b(new_n7144), .O(new_n7168));
  nor2 g06975(.a(new_n7168), .b(new_n7167), .O(new_n7169));
  inv1 g06976(.a(new_n7169), .O(new_n7170));
  nor2 g06977(.a(new_n7170), .b(new_n7131), .O(new_n7171));
  nor2 g06978(.a(new_n7169), .b(new_n7130), .O(new_n7172));
  nor2 g06979(.a(new_n7172), .b(new_n7171), .O(new_n7173));
  inv1 g06980(.a(new_n7173), .O(new_n7174));
  nor2 g06981(.a(new_n6780), .b(new_n6775), .O(new_n7175));
  nor2 g06982(.a(new_n6800), .b(new_n6794), .O(new_n7176));
  inv1 g06983(.a(new_n7176), .O(new_n7177));
  nor2 g06984(.a(new_n6829), .b(new_n6813), .O(new_n7178));
  inv1 g06985(.a(new_n7178), .O(new_n7179));
  nor2 g06986(.a(new_n7179), .b(new_n7177), .O(new_n7180));
  nor2 g06987(.a(new_n7178), .b(new_n7176), .O(new_n7181));
  nor2 g06988(.a(new_n7181), .b(new_n7180), .O(new_n7182));
  nor2 g06989(.a(new_n6856), .b(new_n6850), .O(new_n7183));
  inv1 g06990(.a(new_n7183), .O(new_n7184));
  nor2 g06991(.a(new_n7184), .b(new_n7182), .O(new_n7185));
  inv1 g06992(.a(new_n7182), .O(new_n7186));
  nor2 g06993(.a(new_n7183), .b(new_n7186), .O(new_n7187));
  nor2 g06994(.a(new_n7187), .b(new_n7185), .O(new_n7188));
  nor2 g06995(.a(new_n6836), .b(new_n6806), .O(new_n7189));
  nor2 g06996(.a(new_n6867), .b(new_n6864), .O(new_n7190));
  nor2 g06997(.a(new_n7190), .b(new_n7189), .O(new_n7191));
  inv1 g06998(.a(new_n7189), .O(new_n7192));
  inv1 g06999(.a(new_n7190), .O(new_n7193));
  nor2 g07000(.a(new_n7193), .b(new_n7192), .O(new_n7194));
  nor2 g07001(.a(new_n7194), .b(new_n7191), .O(new_n7195));
  nor2 g07002(.a(new_n7195), .b(new_n7188), .O(new_n7196));
  inv1 g07003(.a(new_n7188), .O(new_n7197));
  inv1 g07004(.a(new_n7195), .O(new_n7198));
  nor2 g07005(.a(new_n7198), .b(new_n7197), .O(new_n7199));
  nor2 g07006(.a(new_n7199), .b(new_n7196), .O(new_n7200));
  inv1 g07007(.a(new_n7200), .O(new_n7201));
  nor2 g07008(.a(new_n7201), .b(new_n7175), .O(new_n7202));
  inv1 g07009(.a(new_n7175), .O(new_n7203));
  nor2 g07010(.a(new_n7200), .b(new_n7203), .O(new_n7204));
  nor2 g07011(.a(new_n7204), .b(new_n7202), .O(new_n7205));
  inv1 g07012(.a(new_n7205), .O(new_n7206));
  nor2 g07013(.a(new_n7206), .b(new_n7174), .O(new_n7207));
  nor2 g07014(.a(new_n7205), .b(new_n7173), .O(new_n7208));
  nor2 g07015(.a(new_n7208), .b(new_n7207), .O(new_n7209));
  inv1 g07016(.a(new_n7209), .O(new_n7210));
  nor2 g07017(.a(new_n7210), .b(new_n7099), .O(new_n7211));
  nor2 g07018(.a(new_n7209), .b(new_n7098), .O(new_n7212));
  nor2 g07019(.a(new_n7212), .b(new_n7211), .O(new_n7213));
  nor2 g07020(.a(new_n6927), .b(new_n6786), .O(new_n7214));
  inv1 g07021(.a(new_n7214), .O(new_n7215));
  nor2 g07022(.a(new_n7215), .b(new_n7213), .O(new_n7216));
  inv1 g07023(.a(new_n7213), .O(new_n7217));
  nor2 g07024(.a(new_n7214), .b(new_n7217), .O(new_n7218));
  nor2 g07025(.a(new_n7218), .b(new_n7216), .O(new_n7219));
  inv1 g07026(.a(new_n7219), .O(new_n7220));
  nor2 g07027(.a(new_n6936), .b(new_n6930), .O(new_n7221));
  nor2 g07028(.a(new_n7221), .b(new_n7220), .O(new_n7222));
  inv1 g07029(.a(new_n7221), .O(new_n7223));
  nor2 g07030(.a(new_n7223), .b(new_n7219), .O(new_n7224));
  nor2 g07031(.a(new_n7224), .b(new_n7222), .O(new_n7225));
  inv1 g07032(.a(new_n7225), .O(\asquared[50] ));
  nor2 g07033(.a(new_n7211), .b(new_n7095), .O(new_n7227));
  inv1 g07034(.a(new_n7227), .O(new_n7228));
  nor2 g07035(.a(new_n7207), .b(new_n7202), .O(new_n7229));
  nor2 g07036(.a(new_n7171), .b(new_n7127), .O(new_n7230));
  nor2 g07037(.a(new_n7199), .b(new_n7191), .O(new_n7231));
  nor2 g07038(.a(new_n7158), .b(new_n7153), .O(new_n7232));
  inv1 g07039(.a(new_n7232), .O(new_n7233));
  nor2 g07040(.a(new_n3533), .b(new_n847), .O(new_n7234));
  nor2 g07041(.a(new_n3722), .b(new_n800), .O(new_n7235));
  nor2 g07042(.a(new_n7235), .b(new_n6964), .O(new_n7236));
  nor2 g07043(.a(new_n5971), .b(new_n800), .O(new_n7237));
  inv1 g07044(.a(new_n7237), .O(new_n7238));
  nor2 g07045(.a(new_n7238), .b(new_n4673), .O(new_n7239));
  nor2 g07046(.a(new_n7239), .b(new_n7236), .O(new_n7240));
  inv1 g07047(.a(new_n7240), .O(new_n7241));
  nor2 g07048(.a(new_n7241), .b(new_n7234), .O(new_n7242));
  inv1 g07049(.a(new_n7234), .O(new_n7243));
  nor2 g07050(.a(new_n7240), .b(new_n7243), .O(new_n7244));
  nor2 g07051(.a(new_n7244), .b(new_n7242), .O(new_n7245));
  nor2 g07052(.a(new_n2433), .b(new_n1493), .O(new_n7246));
  inv1 g07053(.a(new_n7246), .O(new_n7247));
  nor2 g07054(.a(new_n2184), .b(new_n1647), .O(new_n7248));
  nor2 g07055(.a(new_n7248), .b(new_n6949), .O(new_n7249));
  inv1 g07056(.a(new_n7248), .O(new_n7250));
  nor2 g07057(.a(new_n7250), .b(new_n6950), .O(new_n7251));
  nor2 g07058(.a(new_n7251), .b(new_n7249), .O(new_n7252));
  nor2 g07059(.a(new_n7252), .b(new_n7247), .O(new_n7253));
  inv1 g07060(.a(new_n7252), .O(new_n7254));
  nor2 g07061(.a(new_n7254), .b(new_n7246), .O(new_n7255));
  nor2 g07062(.a(new_n7255), .b(new_n7253), .O(new_n7256));
  nor2 g07063(.a(new_n7256), .b(new_n7245), .O(new_n7257));
  inv1 g07064(.a(new_n7245), .O(new_n7258));
  inv1 g07065(.a(new_n7256), .O(new_n7259));
  nor2 g07066(.a(new_n7259), .b(new_n7258), .O(new_n7260));
  nor2 g07067(.a(new_n7260), .b(new_n7257), .O(new_n7261));
  nor2 g07068(.a(new_n7261), .b(new_n7233), .O(new_n7262));
  inv1 g07069(.a(new_n7261), .O(new_n7263));
  nor2 g07070(.a(new_n7263), .b(new_n7232), .O(new_n7264));
  nor2 g07071(.a(new_n7264), .b(new_n7262), .O(new_n7265));
  inv1 g07072(.a(new_n7265), .O(new_n7266));
  nor2 g07073(.a(new_n2826), .b(new_n1199), .O(new_n7267));
  inv1 g07074(.a(new_n7267), .O(new_n7268));
  nor2 g07075(.a(new_n2660), .b(new_n1297), .O(new_n7269));
  nor2 g07076(.a(new_n7269), .b(new_n7010), .O(new_n7270));
  inv1 g07077(.a(new_n7007), .O(new_n7271));
  nor2 g07078(.a(new_n2660), .b(new_n1425), .O(new_n7272));
  inv1 g07079(.a(new_n7272), .O(new_n7273));
  nor2 g07080(.a(new_n7273), .b(new_n7271), .O(new_n7274));
  nor2 g07081(.a(new_n7274), .b(new_n7270), .O(new_n7275));
  nor2 g07082(.a(new_n7275), .b(new_n7268), .O(new_n7276));
  inv1 g07083(.a(new_n7275), .O(new_n7277));
  nor2 g07084(.a(new_n7277), .b(new_n7267), .O(new_n7278));
  nor2 g07085(.a(new_n7278), .b(new_n7276), .O(new_n7279));
  inv1 g07086(.a(new_n7279), .O(new_n7280));
  nor2 g07087(.a(new_n6274), .b(new_n214), .O(new_n7281));
  nor2 g07088(.a(new_n3231), .b(new_n941), .O(new_n7282));
  nor2 g07089(.a(new_n7282), .b(new_n7281), .O(new_n7283));
  inv1 g07090(.a(new_n4097), .O(new_n7284));
  nor2 g07091(.a(new_n6274), .b(new_n941), .O(new_n7285));
  inv1 g07092(.a(new_n7285), .O(new_n7286));
  nor2 g07093(.a(new_n7286), .b(new_n7284), .O(new_n7287));
  nor2 g07094(.a(new_n7287), .b(new_n7283), .O(new_n7288));
  nor2 g07095(.a(new_n7288), .b(new_n7000), .O(new_n7289));
  inv1 g07096(.a(new_n7288), .O(new_n7290));
  nor2 g07097(.a(new_n7290), .b(new_n6999), .O(new_n7291));
  nor2 g07098(.a(new_n7291), .b(new_n7289), .O(new_n7292));
  inv1 g07099(.a(new_n7147), .O(new_n7293));
  inv1 g07100(.a(\a[50] ), .O(new_n7294));
  nor2 g07101(.a(new_n7294), .b(new_n198), .O(new_n7295));
  nor2 g07102(.a(new_n6893), .b(new_n196), .O(new_n7296));
  nor2 g07103(.a(new_n7296), .b(new_n7295), .O(new_n7297));
  nor2 g07104(.a(new_n7294), .b(new_n196), .O(new_n7298));
  inv1 g07105(.a(new_n7298), .O(new_n7299));
  nor2 g07106(.a(new_n7299), .b(new_n6895), .O(new_n7300));
  nor2 g07107(.a(new_n7300), .b(new_n7297), .O(new_n7301));
  nor2 g07108(.a(new_n7301), .b(new_n7293), .O(new_n7302));
  inv1 g07109(.a(new_n7301), .O(new_n7303));
  nor2 g07110(.a(new_n7303), .b(new_n7147), .O(new_n7304));
  nor2 g07111(.a(new_n7304), .b(new_n7302), .O(new_n7305));
  nor2 g07112(.a(new_n7305), .b(new_n7292), .O(new_n7306));
  inv1 g07113(.a(new_n7292), .O(new_n7307));
  inv1 g07114(.a(new_n7305), .O(new_n7308));
  nor2 g07115(.a(new_n7308), .b(new_n7307), .O(new_n7309));
  nor2 g07116(.a(new_n7309), .b(new_n7306), .O(new_n7310));
  nor2 g07117(.a(new_n7310), .b(new_n7280), .O(new_n7311));
  inv1 g07118(.a(new_n7310), .O(new_n7312));
  nor2 g07119(.a(new_n7312), .b(new_n7279), .O(new_n7313));
  nor2 g07120(.a(new_n7313), .b(new_n7311), .O(new_n7314));
  inv1 g07121(.a(new_n7314), .O(new_n7315));
  nor2 g07122(.a(new_n4366), .b(new_n569), .O(new_n7316));
  inv1 g07123(.a(new_n7316), .O(new_n7317));
  nor2 g07124(.a(new_n4682), .b(new_n438), .O(new_n7318));
  nor2 g07125(.a(new_n7318), .b(new_n5907), .O(new_n7319));
  inv1 g07126(.a(new_n6986), .O(new_n7320));
  nor2 g07127(.a(new_n4682), .b(new_n502), .O(new_n7321));
  inv1 g07128(.a(new_n7321), .O(new_n7322));
  nor2 g07129(.a(new_n7322), .b(new_n7320), .O(new_n7323));
  nor2 g07130(.a(new_n7323), .b(new_n7319), .O(new_n7324));
  nor2 g07131(.a(new_n7324), .b(new_n7317), .O(new_n7325));
  inv1 g07132(.a(new_n7324), .O(new_n7326));
  nor2 g07133(.a(new_n7326), .b(new_n7316), .O(new_n7327));
  nor2 g07134(.a(new_n7327), .b(new_n7325), .O(new_n7328));
  inv1 g07135(.a(new_n7328), .O(new_n7329));
  nor2 g07136(.a(new_n4093), .b(new_n613), .O(new_n7330));
  nor2 g07137(.a(new_n4954), .b(new_n363), .O(new_n7331));
  nor2 g07138(.a(new_n7331), .b(new_n7330), .O(new_n7332));
  nor2 g07139(.a(new_n4954), .b(new_n613), .O(new_n7333));
  inv1 g07140(.a(new_n7333), .O(new_n7334));
  nor2 g07141(.a(new_n7334), .b(new_n5991), .O(new_n7335));
  nor2 g07142(.a(new_n7335), .b(new_n7332), .O(new_n7336));
  nor2 g07143(.a(new_n7336), .b(new_n7052), .O(new_n7337));
  inv1 g07144(.a(new_n7336), .O(new_n7338));
  nor2 g07145(.a(new_n7338), .b(new_n7051), .O(new_n7339));
  nor2 g07146(.a(new_n7339), .b(new_n7337), .O(new_n7340));
  nor2 g07147(.a(new_n5796), .b(new_n257), .O(new_n7341));
  inv1 g07148(.a(new_n7341), .O(new_n7342));
  nor2 g07149(.a(new_n5393), .b(new_n295), .O(new_n7343));
  nor2 g07150(.a(new_n3870), .b(new_n699), .O(new_n7344));
  nor2 g07151(.a(new_n7344), .b(new_n7343), .O(new_n7345));
  inv1 g07152(.a(new_n7343), .O(new_n7346));
  inv1 g07153(.a(new_n7344), .O(new_n7347));
  nor2 g07154(.a(new_n7347), .b(new_n7346), .O(new_n7348));
  nor2 g07155(.a(new_n7348), .b(new_n7345), .O(new_n7349));
  nor2 g07156(.a(new_n7349), .b(new_n7342), .O(new_n7350));
  inv1 g07157(.a(new_n7349), .O(new_n7351));
  nor2 g07158(.a(new_n7351), .b(new_n7341), .O(new_n7352));
  nor2 g07159(.a(new_n7352), .b(new_n7350), .O(new_n7353));
  nor2 g07160(.a(new_n7353), .b(new_n7340), .O(new_n7354));
  inv1 g07161(.a(new_n7340), .O(new_n7355));
  inv1 g07162(.a(new_n7353), .O(new_n7356));
  nor2 g07163(.a(new_n7356), .b(new_n7355), .O(new_n7357));
  nor2 g07164(.a(new_n7357), .b(new_n7354), .O(new_n7358));
  nor2 g07165(.a(new_n7358), .b(new_n7329), .O(new_n7359));
  inv1 g07166(.a(new_n7358), .O(new_n7360));
  nor2 g07167(.a(new_n7360), .b(new_n7328), .O(new_n7361));
  nor2 g07168(.a(new_n7361), .b(new_n7359), .O(new_n7362));
  inv1 g07169(.a(new_n7362), .O(new_n7363));
  nor2 g07170(.a(new_n7363), .b(new_n7315), .O(new_n7364));
  nor2 g07171(.a(new_n7362), .b(new_n7314), .O(new_n7365));
  nor2 g07172(.a(new_n7365), .b(new_n7364), .O(new_n7366));
  inv1 g07173(.a(new_n7366), .O(new_n7367));
  nor2 g07174(.a(new_n7367), .b(new_n7266), .O(new_n7368));
  nor2 g07175(.a(new_n7366), .b(new_n7265), .O(new_n7369));
  nor2 g07176(.a(new_n7369), .b(new_n7368), .O(new_n7370));
  inv1 g07177(.a(new_n7370), .O(new_n7371));
  nor2 g07178(.a(new_n7371), .b(new_n7231), .O(new_n7372));
  inv1 g07179(.a(new_n7231), .O(new_n7373));
  nor2 g07180(.a(new_n7370), .b(new_n7373), .O(new_n7374));
  nor2 g07181(.a(new_n7374), .b(new_n7372), .O(new_n7375));
  inv1 g07182(.a(new_n7375), .O(new_n7376));
  nor2 g07183(.a(new_n7376), .b(new_n7230), .O(new_n7377));
  inv1 g07184(.a(new_n7230), .O(new_n7378));
  nor2 g07185(.a(new_n7375), .b(new_n7378), .O(new_n7379));
  nor2 g07186(.a(new_n7379), .b(new_n7377), .O(new_n7380));
  inv1 g07187(.a(new_n7380), .O(new_n7381));
  nor2 g07188(.a(new_n7381), .b(new_n7229), .O(new_n7382));
  inv1 g07189(.a(new_n7229), .O(new_n7383));
  nor2 g07190(.a(new_n7380), .b(new_n7383), .O(new_n7384));
  nor2 g07191(.a(new_n7384), .b(new_n7382), .O(new_n7385));
  inv1 g07192(.a(new_n7385), .O(new_n7386));
  nor2 g07193(.a(new_n7090), .b(new_n7085), .O(new_n7387));
  inv1 g07194(.a(new_n7387), .O(new_n7388));
  nor2 g07195(.a(new_n7123), .b(new_n7117), .O(new_n7389));
  inv1 g07196(.a(new_n7389), .O(new_n7390));
  nor2 g07197(.a(new_n7167), .b(new_n7162), .O(new_n7391));
  inv1 g07198(.a(new_n7391), .O(new_n7392));
  nor2 g07199(.a(new_n7392), .b(new_n7390), .O(new_n7393));
  nor2 g07200(.a(new_n7391), .b(new_n7389), .O(new_n7394));
  nor2 g07201(.a(new_n7394), .b(new_n7393), .O(new_n7395));
  inv1 g07202(.a(new_n7395), .O(new_n7396));
  nor2 g07203(.a(new_n7111), .b(new_n7105), .O(new_n7397));
  inv1 g07204(.a(new_n7397), .O(new_n7398));
  nor2 g07205(.a(new_n7143), .b(new_n7137), .O(new_n7399));
  inv1 g07206(.a(new_n7399), .O(new_n7400));
  nor2 g07207(.a(new_n7400), .b(new_n7398), .O(new_n7401));
  nor2 g07208(.a(new_n7399), .b(new_n7397), .O(new_n7402));
  nor2 g07209(.a(new_n7402), .b(new_n7401), .O(new_n7403));
  inv1 g07210(.a(new_n7403), .O(new_n7404));
  nor2 g07211(.a(new_n6970), .b(new_n6963), .O(new_n7405));
  nor2 g07212(.a(new_n7004), .b(new_n6998), .O(new_n7406));
  nor2 g07213(.a(new_n7406), .b(new_n7405), .O(new_n7407));
  inv1 g07214(.a(new_n7405), .O(new_n7408));
  inv1 g07215(.a(new_n7406), .O(new_n7409));
  nor2 g07216(.a(new_n7409), .b(new_n7408), .O(new_n7410));
  nor2 g07217(.a(new_n7410), .b(new_n7407), .O(new_n7411));
  nor2 g07218(.a(new_n7044), .b(new_n7036), .O(new_n7412));
  nor2 g07219(.a(new_n7412), .b(new_n7411), .O(new_n7413));
  inv1 g07220(.a(new_n7411), .O(new_n7414));
  inv1 g07221(.a(new_n7412), .O(new_n7415));
  nor2 g07222(.a(new_n7415), .b(new_n7414), .O(new_n7416));
  nor2 g07223(.a(new_n7416), .b(new_n7413), .O(new_n7417));
  inv1 g07224(.a(new_n7417), .O(new_n7418));
  nor2 g07225(.a(new_n7418), .b(new_n7404), .O(new_n7419));
  nor2 g07226(.a(new_n7417), .b(new_n7403), .O(new_n7420));
  nor2 g07227(.a(new_n7420), .b(new_n7419), .O(new_n7421));
  inv1 g07228(.a(new_n7421), .O(new_n7422));
  nor2 g07229(.a(new_n7422), .b(new_n7396), .O(new_n7423));
  nor2 g07230(.a(new_n7421), .b(new_n7395), .O(new_n7424));
  nor2 g07231(.a(new_n7424), .b(new_n7423), .O(new_n7425));
  nor2 g07232(.a(new_n7425), .b(new_n7388), .O(new_n7426));
  inv1 g07233(.a(new_n7425), .O(new_n7427));
  nor2 g07234(.a(new_n7427), .b(new_n7387), .O(new_n7428));
  nor2 g07235(.a(new_n7428), .b(new_n7426), .O(new_n7429));
  inv1 g07236(.a(new_n7429), .O(new_n7430));
  nor2 g07237(.a(new_n6978), .b(new_n6972), .O(new_n7431));
  inv1 g07238(.a(new_n7431), .O(new_n7432));
  nor2 g07239(.a(new_n7025), .b(new_n7018), .O(new_n7433));
  inv1 g07240(.a(new_n7433), .O(new_n7434));
  nor2 g07241(.a(new_n7434), .b(new_n7432), .O(new_n7435));
  nor2 g07242(.a(new_n7433), .b(new_n7431), .O(new_n7436));
  nor2 g07243(.a(new_n7436), .b(new_n7435), .O(new_n7437));
  inv1 g07244(.a(new_n7437), .O(new_n7438));
  nor2 g07245(.a(new_n2121), .b(new_n1736), .O(new_n7439));
  nor2 g07246(.a(new_n6958), .b(new_n194), .O(new_n7440));
  nor2 g07247(.a(new_n7440), .b(new_n7439), .O(new_n7441));
  inv1 g07248(.a(new_n7439), .O(new_n7442));
  inv1 g07249(.a(new_n7440), .O(new_n7443));
  nor2 g07250(.a(new_n7443), .b(new_n7442), .O(new_n7444));
  nor2 g07251(.a(new_n7444), .b(new_n7441), .O(new_n7445));
  nor2 g07252(.a(new_n7069), .b(new_n7062), .O(new_n7446));
  nor2 g07253(.a(new_n7446), .b(new_n7445), .O(new_n7447));
  inv1 g07254(.a(new_n7445), .O(new_n7448));
  inv1 g07255(.a(new_n7446), .O(new_n7449));
  nor2 g07256(.a(new_n7449), .b(new_n7448), .O(new_n7450));
  nor2 g07257(.a(new_n7450), .b(new_n7447), .O(new_n7451));
  inv1 g07258(.a(new_n7451), .O(new_n7452));
  nor2 g07259(.a(new_n6994), .b(new_n6987), .O(new_n7453));
  inv1 g07260(.a(new_n7453), .O(new_n7454));
  nor2 g07261(.a(new_n7454), .b(new_n7452), .O(new_n7455));
  nor2 g07262(.a(new_n7453), .b(new_n7451), .O(new_n7456));
  nor2 g07263(.a(new_n7456), .b(new_n7455), .O(new_n7457));
  inv1 g07264(.a(new_n7457), .O(new_n7458));
  nor2 g07265(.a(new_n7458), .b(new_n7438), .O(new_n7459));
  nor2 g07266(.a(new_n7457), .b(new_n7437), .O(new_n7460));
  nor2 g07267(.a(new_n7460), .b(new_n7459), .O(new_n7461));
  inv1 g07268(.a(new_n7461), .O(new_n7462));
  nor2 g07269(.a(new_n7016), .b(new_n7009), .O(new_n7463));
  nor2 g07270(.a(new_n6955), .b(new_n6948), .O(new_n7464));
  nor2 g07271(.a(new_n7464), .b(new_n7463), .O(new_n7465));
  inv1 g07272(.a(new_n7463), .O(new_n7466));
  inv1 g07273(.a(new_n7464), .O(new_n7467));
  nor2 g07274(.a(new_n7467), .b(new_n7466), .O(new_n7468));
  nor2 g07275(.a(new_n7468), .b(new_n7465), .O(new_n7469));
  nor2 g07276(.a(new_n7056), .b(new_n7050), .O(new_n7470));
  nor2 g07277(.a(new_n7470), .b(new_n7469), .O(new_n7471));
  inv1 g07278(.a(new_n7469), .O(new_n7472));
  inv1 g07279(.a(new_n7470), .O(new_n7473));
  nor2 g07280(.a(new_n7473), .b(new_n7472), .O(new_n7474));
  nor2 g07281(.a(new_n7474), .b(new_n7471), .O(new_n7475));
  nor2 g07282(.a(new_n7078), .b(new_n7071), .O(new_n7476));
  inv1 g07283(.a(new_n7476), .O(new_n7477));
  nor2 g07284(.a(new_n7477), .b(new_n7475), .O(new_n7478));
  inv1 g07285(.a(new_n7475), .O(new_n7479));
  nor2 g07286(.a(new_n7476), .b(new_n7479), .O(new_n7480));
  nor2 g07287(.a(new_n7480), .b(new_n7478), .O(new_n7481));
  nor2 g07288(.a(new_n7187), .b(new_n7181), .O(new_n7482));
  inv1 g07289(.a(new_n7482), .O(new_n7483));
  nor2 g07290(.a(new_n7483), .b(new_n7481), .O(new_n7484));
  inv1 g07291(.a(new_n7481), .O(new_n7485));
  nor2 g07292(.a(new_n7482), .b(new_n7485), .O(new_n7486));
  nor2 g07293(.a(new_n7486), .b(new_n7484), .O(new_n7487));
  inv1 g07294(.a(new_n7487), .O(new_n7488));
  nor2 g07295(.a(new_n7081), .b(new_n7028), .O(new_n7489));
  nor2 g07296(.a(new_n7489), .b(new_n7488), .O(new_n7490));
  inv1 g07297(.a(new_n7489), .O(new_n7491));
  nor2 g07298(.a(new_n7491), .b(new_n7487), .O(new_n7492));
  nor2 g07299(.a(new_n7492), .b(new_n7490), .O(new_n7493));
  inv1 g07300(.a(new_n7493), .O(new_n7494));
  nor2 g07301(.a(new_n7494), .b(new_n7462), .O(new_n7495));
  nor2 g07302(.a(new_n7493), .b(new_n7461), .O(new_n7496));
  nor2 g07303(.a(new_n7496), .b(new_n7495), .O(new_n7497));
  inv1 g07304(.a(new_n7497), .O(new_n7498));
  nor2 g07305(.a(new_n7498), .b(new_n7430), .O(new_n7499));
  nor2 g07306(.a(new_n7497), .b(new_n7429), .O(new_n7500));
  nor2 g07307(.a(new_n7500), .b(new_n7499), .O(new_n7501));
  inv1 g07308(.a(new_n7501), .O(new_n7502));
  nor2 g07309(.a(new_n7502), .b(new_n7386), .O(new_n7503));
  nor2 g07310(.a(new_n7501), .b(new_n7385), .O(new_n7504));
  nor2 g07311(.a(new_n7504), .b(new_n7503), .O(new_n7505));
  nor2 g07312(.a(new_n7505), .b(new_n7228), .O(new_n7506));
  inv1 g07313(.a(new_n7505), .O(new_n7507));
  nor2 g07314(.a(new_n7507), .b(new_n7227), .O(new_n7508));
  nor2 g07315(.a(new_n7508), .b(new_n7506), .O(new_n7509));
  inv1 g07316(.a(new_n7509), .O(new_n7510));
  nor2 g07317(.a(new_n7222), .b(new_n7216), .O(new_n7511));
  nor2 g07318(.a(new_n7511), .b(new_n7510), .O(new_n7512));
  inv1 g07319(.a(new_n7511), .O(new_n7513));
  nor2 g07320(.a(new_n7513), .b(new_n7509), .O(new_n7514));
  nor2 g07321(.a(new_n7514), .b(new_n7512), .O(new_n7515));
  inv1 g07322(.a(new_n7515), .O(\asquared[51] ));
  nor2 g07323(.a(new_n7503), .b(new_n7382), .O(new_n7517));
  nor2 g07324(.a(new_n7499), .b(new_n7428), .O(new_n7518));
  nor2 g07325(.a(new_n7495), .b(new_n7490), .O(new_n7519));
  nor2 g07326(.a(new_n7423), .b(new_n7394), .O(new_n7520));
  nor2 g07327(.a(new_n7474), .b(new_n7468), .O(new_n7521));
  inv1 g07328(.a(new_n7521), .O(new_n7522));
  nor2 g07329(.a(new_n3533), .b(new_n941), .O(new_n7523));
  inv1 g07330(.a(new_n7523), .O(new_n7524));
  nor2 g07331(.a(new_n2826), .b(new_n1297), .O(new_n7525));
  nor2 g07332(.a(new_n3057), .b(new_n1199), .O(new_n7526));
  nor2 g07333(.a(new_n7526), .b(new_n7525), .O(new_n7527));
  nor2 g07334(.a(new_n3057), .b(new_n1297), .O(new_n7528));
  inv1 g07335(.a(new_n7528), .O(new_n7529));
  nor2 g07336(.a(new_n7529), .b(new_n7268), .O(new_n7530));
  nor2 g07337(.a(new_n7530), .b(new_n7527), .O(new_n7531));
  nor2 g07338(.a(new_n7531), .b(new_n7524), .O(new_n7532));
  inv1 g07339(.a(new_n7531), .O(new_n7533));
  nor2 g07340(.a(new_n7533), .b(new_n7523), .O(new_n7534));
  nor2 g07341(.a(new_n7534), .b(new_n7532), .O(new_n7535));
  inv1 g07342(.a(new_n7444), .O(new_n7536));
  inv1 g07343(.a(\a[51] ), .O(new_n7537));
  nor2 g07344(.a(new_n7537), .b(new_n198), .O(new_n7538));
  inv1 g07345(.a(new_n7538), .O(new_n7539));
  nor2 g07346(.a(new_n7539), .b(new_n7536), .O(new_n7540));
  nor2 g07347(.a(new_n7538), .b(new_n7444), .O(new_n7541));
  nor2 g07348(.a(new_n7541), .b(new_n7540), .O(new_n7542));
  inv1 g07349(.a(new_n7542), .O(new_n7543));
  nor2 g07350(.a(new_n7294), .b(new_n194), .O(new_n7544));
  inv1 g07351(.a(new_n7544), .O(new_n7545));
  nor2 g07352(.a(new_n7545), .b(new_n2121), .O(new_n7546));
  nor2 g07353(.a(new_n7544), .b(\a[26] ), .O(new_n7547));
  nor2 g07354(.a(new_n7547), .b(new_n7546), .O(new_n7548));
  inv1 g07355(.a(new_n7548), .O(new_n7549));
  nor2 g07356(.a(new_n7549), .b(new_n7543), .O(new_n7550));
  nor2 g07357(.a(new_n7548), .b(new_n7542), .O(new_n7551));
  nor2 g07358(.a(new_n7551), .b(new_n7550), .O(new_n7552));
  inv1 g07359(.a(new_n7552), .O(new_n7553));
  nor2 g07360(.a(new_n7553), .b(new_n7535), .O(new_n7554));
  inv1 g07361(.a(new_n7535), .O(new_n7555));
  nor2 g07362(.a(new_n7552), .b(new_n7555), .O(new_n7556));
  nor2 g07363(.a(new_n7556), .b(new_n7554), .O(new_n7557));
  nor2 g07364(.a(new_n7557), .b(new_n7522), .O(new_n7558));
  inv1 g07365(.a(new_n7557), .O(new_n7559));
  nor2 g07366(.a(new_n7559), .b(new_n7521), .O(new_n7560));
  nor2 g07367(.a(new_n7560), .b(new_n7558), .O(new_n7561));
  inv1 g07368(.a(new_n7561), .O(new_n7562));
  nor2 g07369(.a(new_n2506), .b(new_n1493), .O(new_n7563));
  nor2 g07370(.a(new_n2433), .b(new_n1647), .O(new_n7564));
  nor2 g07371(.a(new_n7564), .b(new_n7563), .O(new_n7565));
  nor2 g07372(.a(new_n2506), .b(new_n1647), .O(new_n7566));
  inv1 g07373(.a(new_n7566), .O(new_n7567));
  nor2 g07374(.a(new_n7567), .b(new_n7247), .O(new_n7568));
  nor2 g07375(.a(new_n7568), .b(new_n7565), .O(new_n7569));
  nor2 g07376(.a(new_n7569), .b(new_n7273), .O(new_n7570));
  inv1 g07377(.a(new_n7569), .O(new_n7571));
  nor2 g07378(.a(new_n7571), .b(new_n7272), .O(new_n7572));
  nor2 g07379(.a(new_n7572), .b(new_n7570), .O(new_n7573));
  nor2 g07380(.a(new_n3231), .b(new_n1086), .O(new_n7574));
  inv1 g07381(.a(new_n7574), .O(new_n7575));
  nor2 g07382(.a(new_n6274), .b(new_n229), .O(new_n7576));
  nor2 g07383(.a(new_n3722), .b(new_n847), .O(new_n7577));
  nor2 g07384(.a(new_n7577), .b(new_n7576), .O(new_n7578));
  inv1 g07385(.a(new_n7576), .O(new_n7579));
  inv1 g07386(.a(new_n7577), .O(new_n7580));
  nor2 g07387(.a(new_n7580), .b(new_n7579), .O(new_n7581));
  nor2 g07388(.a(new_n7581), .b(new_n7578), .O(new_n7582));
  nor2 g07389(.a(new_n7582), .b(new_n7575), .O(new_n7583));
  inv1 g07390(.a(new_n7582), .O(new_n7584));
  nor2 g07391(.a(new_n7584), .b(new_n7574), .O(new_n7585));
  nor2 g07392(.a(new_n7585), .b(new_n7583), .O(new_n7586));
  nor2 g07393(.a(new_n7586), .b(new_n7573), .O(new_n7587));
  inv1 g07394(.a(new_n7573), .O(new_n7588));
  inv1 g07395(.a(new_n7586), .O(new_n7589));
  nor2 g07396(.a(new_n7589), .b(new_n7588), .O(new_n7590));
  nor2 g07397(.a(new_n7590), .b(new_n7587), .O(new_n7591));
  inv1 g07398(.a(new_n7591), .O(new_n7592));
  nor2 g07399(.a(new_n3870), .b(new_n800), .O(new_n7593));
  inv1 g07400(.a(new_n7593), .O(new_n7594));
  nor2 g07401(.a(new_n5971), .b(new_n257), .O(new_n7595));
  nor2 g07402(.a(new_n4093), .b(new_n699), .O(new_n7596));
  nor2 g07403(.a(new_n7596), .b(new_n7595), .O(new_n7597));
  nor2 g07404(.a(new_n5971), .b(new_n699), .O(new_n7598));
  inv1 g07405(.a(new_n7598), .O(new_n7599));
  nor2 g07406(.a(new_n7599), .b(new_n5522), .O(new_n7600));
  nor2 g07407(.a(new_n7600), .b(new_n7597), .O(new_n7601));
  nor2 g07408(.a(new_n7601), .b(new_n7594), .O(new_n7602));
  inv1 g07409(.a(new_n7601), .O(new_n7603));
  nor2 g07410(.a(new_n7603), .b(new_n7593), .O(new_n7604));
  nor2 g07411(.a(new_n7604), .b(new_n7602), .O(new_n7605));
  nor2 g07412(.a(new_n7605), .b(new_n7592), .O(new_n7606));
  inv1 g07413(.a(new_n7605), .O(new_n7607));
  nor2 g07414(.a(new_n7607), .b(new_n7591), .O(new_n7608));
  nor2 g07415(.a(new_n7608), .b(new_n7606), .O(new_n7609));
  inv1 g07416(.a(new_n7609), .O(new_n7610));
  nor2 g07417(.a(new_n2121), .b(new_n1903), .O(new_n7611));
  nor2 g07418(.a(new_n2184), .b(new_n1736), .O(new_n7612));
  nor2 g07419(.a(new_n7612), .b(new_n7611), .O(new_n7613));
  nor2 g07420(.a(new_n2184), .b(new_n1903), .O(new_n7614));
  inv1 g07421(.a(new_n7614), .O(new_n7615));
  nor2 g07422(.a(new_n7615), .b(new_n7442), .O(new_n7616));
  nor2 g07423(.a(new_n7616), .b(new_n7613), .O(new_n7617));
  nor2 g07424(.a(new_n7617), .b(new_n7322), .O(new_n7618));
  inv1 g07425(.a(new_n7617), .O(new_n7619));
  nor2 g07426(.a(new_n7619), .b(new_n7321), .O(new_n7620));
  nor2 g07427(.a(new_n7620), .b(new_n7618), .O(new_n7621));
  nor2 g07428(.a(new_n5796), .b(new_n295), .O(new_n7622));
  nor2 g07429(.a(new_n4366), .b(new_n613), .O(new_n7623));
  nor2 g07430(.a(new_n5393), .b(new_n322), .O(new_n7624));
  nor2 g07431(.a(new_n7624), .b(new_n7623), .O(new_n7625));
  inv1 g07432(.a(new_n6214), .O(new_n7626));
  nor2 g07433(.a(new_n5393), .b(new_n613), .O(new_n7627));
  inv1 g07434(.a(new_n7627), .O(new_n7628));
  nor2 g07435(.a(new_n7628), .b(new_n7626), .O(new_n7629));
  nor2 g07436(.a(new_n7629), .b(new_n7625), .O(new_n7630));
  inv1 g07437(.a(new_n7630), .O(new_n7631));
  nor2 g07438(.a(new_n7631), .b(new_n7622), .O(new_n7632));
  inv1 g07439(.a(new_n7622), .O(new_n7633));
  nor2 g07440(.a(new_n7630), .b(new_n7633), .O(new_n7634));
  nor2 g07441(.a(new_n7634), .b(new_n7632), .O(new_n7635));
  nor2 g07442(.a(new_n5178), .b(new_n363), .O(new_n7636));
  inv1 g07443(.a(new_n7636), .O(new_n7637));
  nor2 g07444(.a(new_n4954), .b(new_n438), .O(new_n7638));
  nor2 g07445(.a(new_n7638), .b(new_n6988), .O(new_n7639));
  nor2 g07446(.a(new_n4954), .b(new_n569), .O(new_n7640));
  inv1 g07447(.a(new_n7640), .O(new_n7641));
  nor2 g07448(.a(new_n7641), .b(new_n7320), .O(new_n7642));
  nor2 g07449(.a(new_n7642), .b(new_n7639), .O(new_n7643));
  nor2 g07450(.a(new_n7643), .b(new_n7637), .O(new_n7644));
  inv1 g07451(.a(new_n7643), .O(new_n7645));
  nor2 g07452(.a(new_n7645), .b(new_n7636), .O(new_n7646));
  nor2 g07453(.a(new_n7646), .b(new_n7644), .O(new_n7647));
  nor2 g07454(.a(new_n7647), .b(new_n7635), .O(new_n7648));
  inv1 g07455(.a(new_n7635), .O(new_n7649));
  inv1 g07456(.a(new_n7647), .O(new_n7650));
  nor2 g07457(.a(new_n7650), .b(new_n7649), .O(new_n7651));
  nor2 g07458(.a(new_n7651), .b(new_n7648), .O(new_n7652));
  inv1 g07459(.a(new_n7652), .O(new_n7653));
  nor2 g07460(.a(new_n7653), .b(new_n7621), .O(new_n7654));
  inv1 g07461(.a(new_n7621), .O(new_n7655));
  nor2 g07462(.a(new_n7652), .b(new_n7655), .O(new_n7656));
  nor2 g07463(.a(new_n7656), .b(new_n7654), .O(new_n7657));
  inv1 g07464(.a(new_n7657), .O(new_n7658));
  nor2 g07465(.a(new_n7658), .b(new_n7610), .O(new_n7659));
  nor2 g07466(.a(new_n7657), .b(new_n7609), .O(new_n7660));
  nor2 g07467(.a(new_n7660), .b(new_n7659), .O(new_n7661));
  inv1 g07468(.a(new_n7661), .O(new_n7662));
  nor2 g07469(.a(new_n7662), .b(new_n7562), .O(new_n7663));
  nor2 g07470(.a(new_n7661), .b(new_n7561), .O(new_n7664));
  nor2 g07471(.a(new_n7664), .b(new_n7663), .O(new_n7665));
  inv1 g07472(.a(new_n7665), .O(new_n7666));
  nor2 g07473(.a(new_n7666), .b(new_n7520), .O(new_n7667));
  inv1 g07474(.a(new_n7520), .O(new_n7668));
  nor2 g07475(.a(new_n7665), .b(new_n7668), .O(new_n7669));
  nor2 g07476(.a(new_n7669), .b(new_n7667), .O(new_n7670));
  inv1 g07477(.a(new_n7670), .O(new_n7671));
  nor2 g07478(.a(new_n7671), .b(new_n7519), .O(new_n7672));
  inv1 g07479(.a(new_n7519), .O(new_n7673));
  nor2 g07480(.a(new_n7670), .b(new_n7673), .O(new_n7674));
  nor2 g07481(.a(new_n7674), .b(new_n7672), .O(new_n7675));
  inv1 g07482(.a(new_n7675), .O(new_n7676));
  nor2 g07483(.a(new_n7676), .b(new_n7518), .O(new_n7677));
  inv1 g07484(.a(new_n7518), .O(new_n7678));
  nor2 g07485(.a(new_n7675), .b(new_n7678), .O(new_n7679));
  nor2 g07486(.a(new_n7679), .b(new_n7677), .O(new_n7680));
  inv1 g07487(.a(new_n7680), .O(new_n7681));
  nor2 g07488(.a(new_n7377), .b(new_n7372), .O(new_n7682));
  nor2 g07489(.a(new_n7486), .b(new_n7480), .O(new_n7683));
  inv1 g07490(.a(new_n7683), .O(new_n7684));
  nor2 g07491(.a(new_n7459), .b(new_n7436), .O(new_n7685));
  inv1 g07492(.a(new_n7685), .O(new_n7686));
  nor2 g07493(.a(new_n7686), .b(new_n7684), .O(new_n7687));
  nor2 g07494(.a(new_n7685), .b(new_n7683), .O(new_n7688));
  nor2 g07495(.a(new_n7688), .b(new_n7687), .O(new_n7689));
  inv1 g07496(.a(new_n7689), .O(new_n7690));
  nor2 g07497(.a(new_n7416), .b(new_n7410), .O(new_n7691));
  inv1 g07498(.a(new_n7691), .O(new_n7692));
  nor2 g07499(.a(new_n7455), .b(new_n7450), .O(new_n7693));
  inv1 g07500(.a(new_n7693), .O(new_n7694));
  nor2 g07501(.a(new_n7694), .b(new_n7692), .O(new_n7695));
  nor2 g07502(.a(new_n7693), .b(new_n7691), .O(new_n7696));
  nor2 g07503(.a(new_n7696), .b(new_n7695), .O(new_n7697));
  nor2 g07504(.a(new_n7313), .b(new_n7306), .O(new_n7698));
  inv1 g07505(.a(new_n7698), .O(new_n7699));
  nor2 g07506(.a(new_n7699), .b(new_n7697), .O(new_n7700));
  inv1 g07507(.a(new_n7697), .O(new_n7701));
  nor2 g07508(.a(new_n7698), .b(new_n7701), .O(new_n7702));
  nor2 g07509(.a(new_n7702), .b(new_n7700), .O(new_n7703));
  inv1 g07510(.a(new_n7703), .O(new_n7704));
  nor2 g07511(.a(new_n7704), .b(new_n7690), .O(new_n7705));
  nor2 g07512(.a(new_n7703), .b(new_n7689), .O(new_n7706));
  nor2 g07513(.a(new_n7706), .b(new_n7705), .O(new_n7707));
  inv1 g07514(.a(new_n7707), .O(new_n7708));
  nor2 g07515(.a(new_n7708), .b(new_n7682), .O(new_n7709));
  inv1 g07516(.a(new_n7682), .O(new_n7710));
  nor2 g07517(.a(new_n7707), .b(new_n7710), .O(new_n7711));
  nor2 g07518(.a(new_n7711), .b(new_n7709), .O(new_n7712));
  inv1 g07519(.a(new_n7712), .O(new_n7713));
  nor2 g07520(.a(new_n7368), .b(new_n7364), .O(new_n7714));
  nor2 g07521(.a(new_n7264), .b(new_n7257), .O(new_n7715));
  inv1 g07522(.a(new_n7715), .O(new_n7716));
  nor2 g07523(.a(new_n7327), .b(new_n7319), .O(new_n7717));
  nor2 g07524(.a(new_n7242), .b(new_n7236), .O(new_n7718));
  nor2 g07525(.a(new_n7718), .b(new_n7717), .O(new_n7719));
  inv1 g07526(.a(new_n7717), .O(new_n7720));
  inv1 g07527(.a(new_n7718), .O(new_n7721));
  nor2 g07528(.a(new_n7721), .b(new_n7720), .O(new_n7722));
  nor2 g07529(.a(new_n7722), .b(new_n7719), .O(new_n7723));
  inv1 g07530(.a(new_n7723), .O(new_n7724));
  nor2 g07531(.a(new_n6958), .b(new_n196), .O(new_n7725));
  inv1 g07532(.a(new_n7725), .O(new_n7726));
  nor2 g07533(.a(new_n6893), .b(new_n203), .O(new_n7727));
  nor2 g07534(.a(new_n6570), .b(new_n214), .O(new_n7728));
  nor2 g07535(.a(new_n7728), .b(new_n7727), .O(new_n7729));
  nor2 g07536(.a(new_n6893), .b(new_n214), .O(new_n7730));
  inv1 g07537(.a(new_n7730), .O(new_n7731));
  nor2 g07538(.a(new_n7731), .b(new_n7000), .O(new_n7732));
  nor2 g07539(.a(new_n7732), .b(new_n7729), .O(new_n7733));
  nor2 g07540(.a(new_n7733), .b(new_n7726), .O(new_n7734));
  inv1 g07541(.a(new_n7733), .O(new_n7735));
  nor2 g07542(.a(new_n7735), .b(new_n7725), .O(new_n7736));
  nor2 g07543(.a(new_n7736), .b(new_n7734), .O(new_n7737));
  nor2 g07544(.a(new_n7737), .b(new_n7724), .O(new_n7738));
  inv1 g07545(.a(new_n7737), .O(new_n7739));
  nor2 g07546(.a(new_n7739), .b(new_n7723), .O(new_n7740));
  nor2 g07547(.a(new_n7740), .b(new_n7738), .O(new_n7741));
  nor2 g07548(.a(new_n7741), .b(new_n7716), .O(new_n7742));
  inv1 g07549(.a(new_n7741), .O(new_n7743));
  nor2 g07550(.a(new_n7743), .b(new_n7715), .O(new_n7744));
  nor2 g07551(.a(new_n7744), .b(new_n7742), .O(new_n7745));
  inv1 g07552(.a(new_n7745), .O(new_n7746));
  nor2 g07553(.a(new_n7419), .b(new_n7402), .O(new_n7747));
  nor2 g07554(.a(new_n7747), .b(new_n7746), .O(new_n7748));
  inv1 g07555(.a(new_n7747), .O(new_n7749));
  nor2 g07556(.a(new_n7749), .b(new_n7745), .O(new_n7750));
  nor2 g07557(.a(new_n7750), .b(new_n7748), .O(new_n7751));
  inv1 g07558(.a(new_n7751), .O(new_n7752));
  nor2 g07559(.a(new_n7752), .b(new_n7714), .O(new_n7753));
  inv1 g07560(.a(new_n7714), .O(new_n7754));
  nor2 g07561(.a(new_n7751), .b(new_n7754), .O(new_n7755));
  nor2 g07562(.a(new_n7755), .b(new_n7753), .O(new_n7756));
  inv1 g07563(.a(new_n7756), .O(new_n7757));
  nor2 g07564(.a(new_n7352), .b(new_n7345), .O(new_n7758));
  nor2 g07565(.a(new_n7339), .b(new_n7332), .O(new_n7759));
  nor2 g07566(.a(new_n7759), .b(new_n7758), .O(new_n7760));
  inv1 g07567(.a(new_n7758), .O(new_n7761));
  inv1 g07568(.a(new_n7759), .O(new_n7762));
  nor2 g07569(.a(new_n7762), .b(new_n7761), .O(new_n7763));
  nor2 g07570(.a(new_n7763), .b(new_n7760), .O(new_n7764));
  nor2 g07571(.a(new_n7255), .b(new_n7249), .O(new_n7765));
  nor2 g07572(.a(new_n7765), .b(new_n7764), .O(new_n7766));
  inv1 g07573(.a(new_n7764), .O(new_n7767));
  inv1 g07574(.a(new_n7765), .O(new_n7768));
  nor2 g07575(.a(new_n7768), .b(new_n7767), .O(new_n7769));
  nor2 g07576(.a(new_n7769), .b(new_n7766), .O(new_n7770));
  nor2 g07577(.a(new_n7361), .b(new_n7354), .O(new_n7771));
  inv1 g07578(.a(new_n7771), .O(new_n7772));
  nor2 g07579(.a(new_n7772), .b(new_n7770), .O(new_n7773));
  inv1 g07580(.a(new_n7770), .O(new_n7774));
  nor2 g07581(.a(new_n7771), .b(new_n7774), .O(new_n7775));
  nor2 g07582(.a(new_n7775), .b(new_n7773), .O(new_n7776));
  inv1 g07583(.a(new_n7776), .O(new_n7777));
  nor2 g07584(.a(new_n7291), .b(new_n7283), .O(new_n7778));
  nor2 g07585(.a(new_n7278), .b(new_n7270), .O(new_n7779));
  nor2 g07586(.a(new_n7779), .b(new_n7778), .O(new_n7780));
  inv1 g07587(.a(new_n7778), .O(new_n7781));
  inv1 g07588(.a(new_n7779), .O(new_n7782));
  nor2 g07589(.a(new_n7782), .b(new_n7781), .O(new_n7783));
  nor2 g07590(.a(new_n7783), .b(new_n7780), .O(new_n7784));
  nor2 g07591(.a(new_n7304), .b(new_n7297), .O(new_n7785));
  nor2 g07592(.a(new_n7785), .b(new_n7784), .O(new_n7786));
  inv1 g07593(.a(new_n7784), .O(new_n7787));
  inv1 g07594(.a(new_n7785), .O(new_n7788));
  nor2 g07595(.a(new_n7788), .b(new_n7787), .O(new_n7789));
  nor2 g07596(.a(new_n7789), .b(new_n7786), .O(new_n7790));
  inv1 g07597(.a(new_n7790), .O(new_n7791));
  nor2 g07598(.a(new_n7791), .b(new_n7777), .O(new_n7792));
  nor2 g07599(.a(new_n7790), .b(new_n7776), .O(new_n7793));
  nor2 g07600(.a(new_n7793), .b(new_n7792), .O(new_n7794));
  inv1 g07601(.a(new_n7794), .O(new_n7795));
  nor2 g07602(.a(new_n7795), .b(new_n7757), .O(new_n7796));
  nor2 g07603(.a(new_n7794), .b(new_n7756), .O(new_n7797));
  nor2 g07604(.a(new_n7797), .b(new_n7796), .O(new_n7798));
  inv1 g07605(.a(new_n7798), .O(new_n7799));
  nor2 g07606(.a(new_n7799), .b(new_n7713), .O(new_n7800));
  nor2 g07607(.a(new_n7798), .b(new_n7712), .O(new_n7801));
  nor2 g07608(.a(new_n7801), .b(new_n7800), .O(new_n7802));
  inv1 g07609(.a(new_n7802), .O(new_n7803));
  nor2 g07610(.a(new_n7803), .b(new_n7681), .O(new_n7804));
  nor2 g07611(.a(new_n7802), .b(new_n7680), .O(new_n7805));
  nor2 g07612(.a(new_n7805), .b(new_n7804), .O(new_n7806));
  inv1 g07613(.a(new_n7806), .O(new_n7807));
  nor2 g07614(.a(new_n7807), .b(new_n7517), .O(new_n7808));
  inv1 g07615(.a(new_n7517), .O(new_n7809));
  nor2 g07616(.a(new_n7806), .b(new_n7809), .O(new_n7810));
  nor2 g07617(.a(new_n7810), .b(new_n7808), .O(new_n7811));
  inv1 g07618(.a(new_n7811), .O(new_n7812));
  nor2 g07619(.a(new_n7512), .b(new_n7506), .O(new_n7813));
  nor2 g07620(.a(new_n7813), .b(new_n7812), .O(new_n7814));
  inv1 g07621(.a(new_n7813), .O(new_n7815));
  nor2 g07622(.a(new_n7815), .b(new_n7811), .O(new_n7816));
  nor2 g07623(.a(new_n7816), .b(new_n7814), .O(new_n7817));
  inv1 g07624(.a(new_n7817), .O(\asquared[52] ));
  nor2 g07625(.a(new_n7804), .b(new_n7677), .O(new_n7819));
  inv1 g07626(.a(new_n7819), .O(new_n7820));
  nor2 g07627(.a(new_n7796), .b(new_n7753), .O(new_n7821));
  inv1 g07628(.a(new_n7821), .O(new_n7822));
  nor2 g07629(.a(new_n7705), .b(new_n7688), .O(new_n7823));
  nor2 g07630(.a(new_n7792), .b(new_n7775), .O(new_n7824));
  nor2 g07631(.a(new_n4093), .b(new_n800), .O(new_n7825));
  inv1 g07632(.a(new_n7825), .O(new_n7826));
  nor2 g07633(.a(new_n5971), .b(new_n295), .O(new_n7827));
  nor2 g07634(.a(new_n5796), .b(new_n322), .O(new_n7828));
  nor2 g07635(.a(new_n7828), .b(new_n7827), .O(new_n7829));
  nor2 g07636(.a(new_n5971), .b(new_n322), .O(new_n7830));
  inv1 g07637(.a(new_n7830), .O(new_n7831));
  nor2 g07638(.a(new_n7831), .b(new_n7633), .O(new_n7832));
  nor2 g07639(.a(new_n7832), .b(new_n7829), .O(new_n7833));
  nor2 g07640(.a(new_n7833), .b(new_n7826), .O(new_n7834));
  inv1 g07641(.a(new_n7833), .O(new_n7835));
  nor2 g07642(.a(new_n7835), .b(new_n7825), .O(new_n7836));
  nor2 g07643(.a(new_n7836), .b(new_n7834), .O(new_n7837));
  nor2 g07644(.a(new_n5178), .b(new_n438), .O(new_n7838));
  inv1 g07645(.a(new_n7838), .O(new_n7839));
  nor2 g07646(.a(new_n4954), .b(new_n502), .O(new_n7840));
  nor2 g07647(.a(new_n7840), .b(new_n6450), .O(new_n7841));
  nor2 g07648(.a(new_n7641), .b(new_n7322), .O(new_n7842));
  nor2 g07649(.a(new_n7842), .b(new_n7841), .O(new_n7843));
  nor2 g07650(.a(new_n7843), .b(new_n7839), .O(new_n7844));
  inv1 g07651(.a(new_n7843), .O(new_n7845));
  nor2 g07652(.a(new_n7845), .b(new_n7838), .O(new_n7846));
  nor2 g07653(.a(new_n7846), .b(new_n7844), .O(new_n7847));
  nor2 g07654(.a(new_n6570), .b(new_n229), .O(new_n7848));
  inv1 g07655(.a(new_n7848), .O(new_n7849));
  nor2 g07656(.a(new_n3870), .b(new_n847), .O(new_n7850));
  nor2 g07657(.a(new_n6274), .b(new_n257), .O(new_n7851));
  nor2 g07658(.a(new_n7851), .b(new_n7850), .O(new_n7852));
  nor2 g07659(.a(new_n6274), .b(new_n847), .O(new_n7853));
  inv1 g07660(.a(new_n7853), .O(new_n7854));
  nor2 g07661(.a(new_n7854), .b(new_n5259), .O(new_n7855));
  nor2 g07662(.a(new_n7855), .b(new_n7852), .O(new_n7856));
  nor2 g07663(.a(new_n7856), .b(new_n7849), .O(new_n7857));
  inv1 g07664(.a(new_n7856), .O(new_n7858));
  nor2 g07665(.a(new_n7858), .b(new_n7848), .O(new_n7859));
  nor2 g07666(.a(new_n7859), .b(new_n7857), .O(new_n7860));
  nor2 g07667(.a(new_n7860), .b(new_n7847), .O(new_n7861));
  inv1 g07668(.a(new_n7847), .O(new_n7862));
  inv1 g07669(.a(new_n7860), .O(new_n7863));
  nor2 g07670(.a(new_n7863), .b(new_n7862), .O(new_n7864));
  nor2 g07671(.a(new_n7864), .b(new_n7861), .O(new_n7865));
  inv1 g07672(.a(new_n7865), .O(new_n7866));
  nor2 g07673(.a(new_n7866), .b(new_n7837), .O(new_n7867));
  inv1 g07674(.a(new_n7837), .O(new_n7868));
  nor2 g07675(.a(new_n7865), .b(new_n7868), .O(new_n7869));
  nor2 g07676(.a(new_n7869), .b(new_n7867), .O(new_n7870));
  nor2 g07677(.a(new_n3533), .b(new_n1086), .O(new_n7871));
  nor2 g07678(.a(new_n2826), .b(new_n1425), .O(new_n7872));
  nor2 g07679(.a(new_n7872), .b(new_n7528), .O(new_n7873));
  inv1 g07680(.a(new_n7525), .O(new_n7874));
  nor2 g07681(.a(new_n3057), .b(new_n1425), .O(new_n7875));
  inv1 g07682(.a(new_n7875), .O(new_n7876));
  nor2 g07683(.a(new_n7876), .b(new_n7874), .O(new_n7877));
  nor2 g07684(.a(new_n7877), .b(new_n7873), .O(new_n7878));
  inv1 g07685(.a(new_n7878), .O(new_n7879));
  nor2 g07686(.a(new_n7879), .b(new_n7871), .O(new_n7880));
  inv1 g07687(.a(new_n7871), .O(new_n7881));
  nor2 g07688(.a(new_n7878), .b(new_n7881), .O(new_n7882));
  nor2 g07689(.a(new_n7882), .b(new_n7880), .O(new_n7883));
  nor2 g07690(.a(new_n2660), .b(new_n1493), .O(new_n7884));
  inv1 g07691(.a(new_n7884), .O(new_n7885));
  nor2 g07692(.a(new_n2433), .b(new_n1736), .O(new_n7886));
  nor2 g07693(.a(new_n7886), .b(new_n7566), .O(new_n7887));
  inv1 g07694(.a(new_n7564), .O(new_n7888));
  nor2 g07695(.a(new_n2506), .b(new_n1736), .O(new_n7889));
  inv1 g07696(.a(new_n7889), .O(new_n7890));
  nor2 g07697(.a(new_n7890), .b(new_n7888), .O(new_n7891));
  nor2 g07698(.a(new_n7891), .b(new_n7887), .O(new_n7892));
  nor2 g07699(.a(new_n7892), .b(new_n7885), .O(new_n7893));
  inv1 g07700(.a(new_n7892), .O(new_n7894));
  nor2 g07701(.a(new_n7894), .b(new_n7884), .O(new_n7895));
  nor2 g07702(.a(new_n7895), .b(new_n7893), .O(new_n7896));
  nor2 g07703(.a(new_n7896), .b(new_n7883), .O(new_n7897));
  inv1 g07704(.a(new_n7883), .O(new_n7898));
  inv1 g07705(.a(new_n7896), .O(new_n7899));
  nor2 g07706(.a(new_n7899), .b(new_n7898), .O(new_n7900));
  nor2 g07707(.a(new_n7900), .b(new_n7897), .O(new_n7901));
  inv1 g07708(.a(new_n7901), .O(new_n7902));
  nor2 g07709(.a(new_n5393), .b(new_n363), .O(new_n7903));
  nor2 g07710(.a(new_n4425), .b(new_n613), .O(new_n7904));
  nor2 g07711(.a(new_n7904), .b(new_n7903), .O(new_n7905));
  nor2 g07712(.a(new_n7628), .b(new_n6677), .O(new_n7906));
  nor2 g07713(.a(new_n7906), .b(new_n7905), .O(new_n7907));
  nor2 g07714(.a(new_n7907), .b(new_n5293), .O(new_n7908));
  inv1 g07715(.a(new_n7907), .O(new_n7909));
  nor2 g07716(.a(new_n7909), .b(new_n5292), .O(new_n7910));
  nor2 g07717(.a(new_n7910), .b(new_n7908), .O(new_n7911));
  nor2 g07718(.a(new_n7911), .b(new_n7902), .O(new_n7912));
  inv1 g07719(.a(new_n7911), .O(new_n7913));
  nor2 g07720(.a(new_n7913), .b(new_n7901), .O(new_n7914));
  nor2 g07721(.a(new_n7914), .b(new_n7912), .O(new_n7915));
  nor2 g07722(.a(new_n7915), .b(new_n7870), .O(new_n7916));
  inv1 g07723(.a(new_n7870), .O(new_n7917));
  inv1 g07724(.a(new_n7915), .O(new_n7918));
  nor2 g07725(.a(new_n7918), .b(new_n7917), .O(new_n7919));
  nor2 g07726(.a(new_n7919), .b(new_n7916), .O(new_n7920));
  inv1 g07727(.a(new_n7920), .O(new_n7921));
  nor2 g07728(.a(new_n7921), .b(new_n7824), .O(new_n7922));
  inv1 g07729(.a(new_n7824), .O(new_n7923));
  nor2 g07730(.a(new_n7920), .b(new_n7923), .O(new_n7924));
  nor2 g07731(.a(new_n7924), .b(new_n7922), .O(new_n7925));
  inv1 g07732(.a(new_n7925), .O(new_n7926));
  nor2 g07733(.a(new_n7926), .b(new_n7823), .O(new_n7927));
  inv1 g07734(.a(new_n7823), .O(new_n7928));
  nor2 g07735(.a(new_n7925), .b(new_n7928), .O(new_n7929));
  nor2 g07736(.a(new_n7929), .b(new_n7927), .O(new_n7930));
  nor2 g07737(.a(new_n7930), .b(new_n7822), .O(new_n7931));
  inv1 g07738(.a(new_n7930), .O(new_n7932));
  nor2 g07739(.a(new_n7932), .b(new_n7821), .O(new_n7933));
  nor2 g07740(.a(new_n7933), .b(new_n7931), .O(new_n7934));
  inv1 g07741(.a(new_n7934), .O(new_n7935));
  nor2 g07742(.a(new_n7800), .b(new_n7709), .O(new_n7936));
  nor2 g07743(.a(new_n7936), .b(new_n7935), .O(new_n7937));
  inv1 g07744(.a(new_n7936), .O(new_n7938));
  nor2 g07745(.a(new_n7938), .b(new_n7934), .O(new_n7939));
  nor2 g07746(.a(new_n7939), .b(new_n7937), .O(new_n7940));
  inv1 g07747(.a(new_n7940), .O(new_n7941));
  nor2 g07748(.a(new_n7672), .b(new_n7667), .O(new_n7942));
  inv1 g07749(.a(new_n7942), .O(new_n7943));
  nor2 g07750(.a(new_n7769), .b(new_n7763), .O(new_n7944));
  inv1 g07751(.a(new_n7944), .O(new_n7945));
  nor2 g07752(.a(new_n7789), .b(new_n7783), .O(new_n7946));
  nor2 g07753(.a(new_n3231), .b(new_n1199), .O(new_n7947));
  inv1 g07754(.a(new_n7947), .O(new_n7948));
  nor2 g07755(.a(new_n6958), .b(new_n203), .O(new_n7949));
  nor2 g07756(.a(new_n7949), .b(new_n7298), .O(new_n7950));
  nor2 g07757(.a(new_n7294), .b(new_n203), .O(new_n7951));
  inv1 g07758(.a(new_n7951), .O(new_n7952));
  nor2 g07759(.a(new_n7952), .b(new_n7726), .O(new_n7953));
  nor2 g07760(.a(new_n7953), .b(new_n7950), .O(new_n7954));
  nor2 g07761(.a(new_n7954), .b(new_n7948), .O(new_n7955));
  inv1 g07762(.a(new_n7954), .O(new_n7956));
  nor2 g07763(.a(new_n7956), .b(new_n7947), .O(new_n7957));
  nor2 g07764(.a(new_n7957), .b(new_n7955), .O(new_n7958));
  nor2 g07765(.a(new_n7958), .b(new_n7946), .O(new_n7959));
  inv1 g07766(.a(new_n7946), .O(new_n7960));
  inv1 g07767(.a(new_n7958), .O(new_n7961));
  nor2 g07768(.a(new_n7961), .b(new_n7960), .O(new_n7962));
  nor2 g07769(.a(new_n7962), .b(new_n7959), .O(new_n7963));
  nor2 g07770(.a(new_n7963), .b(new_n7945), .O(new_n7964));
  inv1 g07771(.a(new_n7963), .O(new_n7965));
  nor2 g07772(.a(new_n7965), .b(new_n7944), .O(new_n7966));
  nor2 g07773(.a(new_n7966), .b(new_n7964), .O(new_n7967));
  nor2 g07774(.a(new_n7748), .b(new_n7744), .O(new_n7968));
  inv1 g07775(.a(new_n7968), .O(new_n7969));
  nor2 g07776(.a(new_n7969), .b(new_n7967), .O(new_n7970));
  inv1 g07777(.a(new_n7967), .O(new_n7971));
  nor2 g07778(.a(new_n7968), .b(new_n7971), .O(new_n7972));
  nor2 g07779(.a(new_n7972), .b(new_n7970), .O(new_n7973));
  inv1 g07780(.a(new_n7973), .O(new_n7974));
  nor2 g07781(.a(new_n7654), .b(new_n7648), .O(new_n7975));
  inv1 g07782(.a(new_n7546), .O(new_n7976));
  nor2 g07783(.a(new_n7537), .b(new_n194), .O(new_n7977));
  nor2 g07784(.a(new_n7977), .b(new_n7614), .O(new_n7978));
  inv1 g07785(.a(new_n7977), .O(new_n7979));
  nor2 g07786(.a(new_n7979), .b(new_n7615), .O(new_n7980));
  nor2 g07787(.a(new_n7980), .b(new_n7978), .O(new_n7981));
  inv1 g07788(.a(new_n7981), .O(new_n7982));
  nor2 g07789(.a(new_n7982), .b(new_n7976), .O(new_n7983));
  nor2 g07790(.a(new_n7981), .b(new_n7546), .O(new_n7984));
  nor2 g07791(.a(new_n7984), .b(new_n7983), .O(new_n7985));
  inv1 g07792(.a(new_n7985), .O(new_n7986));
  nor2 g07793(.a(new_n7620), .b(new_n7613), .O(new_n7987));
  inv1 g07794(.a(new_n7987), .O(new_n7988));
  nor2 g07795(.a(new_n7988), .b(new_n7986), .O(new_n7989));
  nor2 g07796(.a(new_n7987), .b(new_n7985), .O(new_n7990));
  nor2 g07797(.a(new_n7990), .b(new_n7989), .O(new_n7991));
  inv1 g07798(.a(new_n7991), .O(new_n7992));
  nor2 g07799(.a(new_n7738), .b(new_n7722), .O(new_n7993));
  nor2 g07800(.a(new_n7993), .b(new_n7992), .O(new_n7994));
  inv1 g07801(.a(new_n7993), .O(new_n7995));
  nor2 g07802(.a(new_n7995), .b(new_n7991), .O(new_n7996));
  nor2 g07803(.a(new_n7996), .b(new_n7994), .O(new_n7997));
  inv1 g07804(.a(new_n7997), .O(new_n7998));
  nor2 g07805(.a(new_n7998), .b(new_n7975), .O(new_n7999));
  inv1 g07806(.a(new_n7975), .O(new_n8000));
  nor2 g07807(.a(new_n7997), .b(new_n8000), .O(new_n8001));
  nor2 g07808(.a(new_n8001), .b(new_n7999), .O(new_n8002));
  inv1 g07809(.a(new_n8002), .O(new_n8003));
  nor2 g07810(.a(new_n8003), .b(new_n7974), .O(new_n8004));
  nor2 g07811(.a(new_n8002), .b(new_n7973), .O(new_n8005));
  nor2 g07812(.a(new_n8005), .b(new_n8004), .O(new_n8006));
  nor2 g07813(.a(new_n8006), .b(new_n7943), .O(new_n8007));
  inv1 g07814(.a(new_n8006), .O(new_n8008));
  nor2 g07815(.a(new_n8008), .b(new_n7942), .O(new_n8009));
  nor2 g07816(.a(new_n8009), .b(new_n8007), .O(new_n8010));
  inv1 g07817(.a(new_n8010), .O(new_n8011));
  nor2 g07818(.a(new_n7560), .b(new_n7554), .O(new_n8012));
  inv1 g07819(.a(new_n8012), .O(new_n8013));
  nor2 g07820(.a(new_n7550), .b(new_n7540), .O(new_n8014));
  inv1 g07821(.a(new_n8014), .O(new_n8015));
  nor2 g07822(.a(new_n7646), .b(new_n7639), .O(new_n8016));
  nor2 g07823(.a(new_n8016), .b(new_n8015), .O(new_n8017));
  inv1 g07824(.a(new_n8016), .O(new_n8018));
  nor2 g07825(.a(new_n8018), .b(new_n8014), .O(new_n8019));
  nor2 g07826(.a(new_n8019), .b(new_n8017), .O(new_n8020));
  nor2 g07827(.a(new_n3722), .b(new_n941), .O(new_n8021));
  nor2 g07828(.a(new_n8021), .b(new_n7730), .O(new_n8022));
  inv1 g07829(.a(new_n8021), .O(new_n8023));
  nor2 g07830(.a(new_n8023), .b(new_n7731), .O(new_n8024));
  nor2 g07831(.a(new_n8024), .b(new_n8022), .O(new_n8025));
  inv1 g07832(.a(\a[52] ), .O(new_n8026));
  nor2 g07833(.a(new_n8026), .b(new_n198), .O(new_n8027));
  inv1 g07834(.a(new_n8027), .O(new_n8028));
  nor2 g07835(.a(new_n8028), .b(new_n8025), .O(new_n8029));
  inv1 g07836(.a(new_n8025), .O(new_n8030));
  nor2 g07837(.a(new_n8027), .b(new_n8030), .O(new_n8031));
  nor2 g07838(.a(new_n8031), .b(new_n8029), .O(new_n8032));
  inv1 g07839(.a(new_n8032), .O(new_n8033));
  nor2 g07840(.a(new_n8033), .b(new_n8020), .O(new_n8034));
  inv1 g07841(.a(new_n8020), .O(new_n8035));
  nor2 g07842(.a(new_n8032), .b(new_n8035), .O(new_n8036));
  nor2 g07843(.a(new_n8036), .b(new_n8034), .O(new_n8037));
  nor2 g07844(.a(new_n8037), .b(new_n8013), .O(new_n8038));
  inv1 g07845(.a(new_n8037), .O(new_n8039));
  nor2 g07846(.a(new_n8039), .b(new_n8012), .O(new_n8040));
  nor2 g07847(.a(new_n8040), .b(new_n8038), .O(new_n8041));
  nor2 g07848(.a(new_n7702), .b(new_n7696), .O(new_n8042));
  inv1 g07849(.a(new_n8042), .O(new_n8043));
  nor2 g07850(.a(new_n8043), .b(new_n8041), .O(new_n8044));
  inv1 g07851(.a(new_n8041), .O(new_n8045));
  nor2 g07852(.a(new_n8042), .b(new_n8045), .O(new_n8046));
  nor2 g07853(.a(new_n8046), .b(new_n8044), .O(new_n8047));
  inv1 g07854(.a(new_n8047), .O(new_n8048));
  nor2 g07855(.a(new_n7663), .b(new_n7659), .O(new_n8049));
  nor2 g07856(.a(new_n7585), .b(new_n7578), .O(new_n8050));
  nor2 g07857(.a(new_n7632), .b(new_n7625), .O(new_n8051));
  nor2 g07858(.a(new_n8051), .b(new_n8050), .O(new_n8052));
  inv1 g07859(.a(new_n8050), .O(new_n8053));
  inv1 g07860(.a(new_n8051), .O(new_n8054));
  nor2 g07861(.a(new_n8054), .b(new_n8053), .O(new_n8055));
  nor2 g07862(.a(new_n8055), .b(new_n8052), .O(new_n8056));
  nor2 g07863(.a(new_n7572), .b(new_n7565), .O(new_n8057));
  nor2 g07864(.a(new_n8057), .b(new_n8056), .O(new_n8058));
  inv1 g07865(.a(new_n8056), .O(new_n8059));
  inv1 g07866(.a(new_n8057), .O(new_n8060));
  nor2 g07867(.a(new_n8060), .b(new_n8059), .O(new_n8061));
  nor2 g07868(.a(new_n8061), .b(new_n8058), .O(new_n8062));
  inv1 g07869(.a(new_n8062), .O(new_n8063));
  nor2 g07870(.a(new_n7534), .b(new_n7527), .O(new_n8064));
  nor2 g07871(.a(new_n7736), .b(new_n7729), .O(new_n8065));
  nor2 g07872(.a(new_n8065), .b(new_n8064), .O(new_n8066));
  inv1 g07873(.a(new_n8064), .O(new_n8067));
  inv1 g07874(.a(new_n8065), .O(new_n8068));
  nor2 g07875(.a(new_n8068), .b(new_n8067), .O(new_n8069));
  nor2 g07876(.a(new_n8069), .b(new_n8066), .O(new_n8070));
  nor2 g07877(.a(new_n7604), .b(new_n7597), .O(new_n8071));
  nor2 g07878(.a(new_n8071), .b(new_n8070), .O(new_n8072));
  inv1 g07879(.a(new_n8070), .O(new_n8073));
  inv1 g07880(.a(new_n8071), .O(new_n8074));
  nor2 g07881(.a(new_n8074), .b(new_n8073), .O(new_n8075));
  nor2 g07882(.a(new_n8075), .b(new_n8072), .O(new_n8076));
  nor2 g07883(.a(new_n7606), .b(new_n7587), .O(new_n8077));
  inv1 g07884(.a(new_n8077), .O(new_n8078));
  nor2 g07885(.a(new_n8078), .b(new_n8076), .O(new_n8079));
  inv1 g07886(.a(new_n8076), .O(new_n8080));
  nor2 g07887(.a(new_n8077), .b(new_n8080), .O(new_n8081));
  nor2 g07888(.a(new_n8081), .b(new_n8079), .O(new_n8082));
  inv1 g07889(.a(new_n8082), .O(new_n8083));
  nor2 g07890(.a(new_n8083), .b(new_n8063), .O(new_n8084));
  nor2 g07891(.a(new_n8082), .b(new_n8062), .O(new_n8085));
  nor2 g07892(.a(new_n8085), .b(new_n8084), .O(new_n8086));
  inv1 g07893(.a(new_n8086), .O(new_n8087));
  nor2 g07894(.a(new_n8087), .b(new_n8049), .O(new_n8088));
  inv1 g07895(.a(new_n8049), .O(new_n8089));
  nor2 g07896(.a(new_n8086), .b(new_n8089), .O(new_n8090));
  nor2 g07897(.a(new_n8090), .b(new_n8088), .O(new_n8091));
  inv1 g07898(.a(new_n8091), .O(new_n8092));
  nor2 g07899(.a(new_n8092), .b(new_n8048), .O(new_n8093));
  nor2 g07900(.a(new_n8091), .b(new_n8047), .O(new_n8094));
  nor2 g07901(.a(new_n8094), .b(new_n8093), .O(new_n8095));
  inv1 g07902(.a(new_n8095), .O(new_n8096));
  nor2 g07903(.a(new_n8096), .b(new_n8011), .O(new_n8097));
  nor2 g07904(.a(new_n8095), .b(new_n8010), .O(new_n8098));
  nor2 g07905(.a(new_n8098), .b(new_n8097), .O(new_n8099));
  inv1 g07906(.a(new_n8099), .O(new_n8100));
  nor2 g07907(.a(new_n8100), .b(new_n7941), .O(new_n8101));
  nor2 g07908(.a(new_n8099), .b(new_n7940), .O(new_n8102));
  nor2 g07909(.a(new_n8102), .b(new_n8101), .O(new_n8103));
  nor2 g07910(.a(new_n8103), .b(new_n7820), .O(new_n8104));
  inv1 g07911(.a(new_n8103), .O(new_n8105));
  nor2 g07912(.a(new_n8105), .b(new_n7819), .O(new_n8106));
  nor2 g07913(.a(new_n8106), .b(new_n8104), .O(new_n8107));
  nor2 g07914(.a(new_n7814), .b(new_n7810), .O(new_n8108));
  inv1 g07915(.a(new_n8108), .O(new_n8109));
  nor2 g07916(.a(new_n8109), .b(new_n8107), .O(new_n8110));
  inv1 g07917(.a(new_n8107), .O(new_n8111));
  nor2 g07918(.a(new_n8108), .b(new_n8111), .O(new_n8112));
  nor2 g07919(.a(new_n8112), .b(new_n8110), .O(new_n8113));
  inv1 g07920(.a(new_n8113), .O(\asquared[53] ));
  nor2 g07921(.a(new_n8101), .b(new_n7937), .O(new_n8115));
  nor2 g07922(.a(new_n8097), .b(new_n8009), .O(new_n8116));
  nor2 g07923(.a(new_n8093), .b(new_n8088), .O(new_n8117));
  nor2 g07924(.a(new_n7966), .b(new_n7959), .O(new_n8118));
  inv1 g07925(.a(new_n8118), .O(new_n8119));
  nor2 g07926(.a(new_n3533), .b(new_n1199), .O(new_n8120));
  inv1 g07927(.a(new_n8120), .O(new_n8121));
  nor2 g07928(.a(new_n3231), .b(new_n1297), .O(new_n8122));
  nor2 g07929(.a(new_n8122), .b(new_n7875), .O(new_n8123));
  nor2 g07930(.a(new_n3231), .b(new_n1425), .O(new_n8124));
  inv1 g07931(.a(new_n8124), .O(new_n8125));
  nor2 g07932(.a(new_n8125), .b(new_n7529), .O(new_n8126));
  nor2 g07933(.a(new_n8126), .b(new_n8123), .O(new_n8127));
  nor2 g07934(.a(new_n8127), .b(new_n8121), .O(new_n8128));
  inv1 g07935(.a(new_n8127), .O(new_n8129));
  nor2 g07936(.a(new_n8129), .b(new_n8120), .O(new_n8130));
  nor2 g07937(.a(new_n8130), .b(new_n8128), .O(new_n8131));
  inv1 g07938(.a(new_n8131), .O(new_n8132));
  nor2 g07939(.a(new_n7537), .b(new_n196), .O(new_n8133));
  nor2 g07940(.a(new_n8133), .b(new_n7951), .O(new_n8134));
  nor2 g07941(.a(new_n7537), .b(new_n203), .O(new_n8135));
  inv1 g07942(.a(new_n8135), .O(new_n8136));
  nor2 g07943(.a(new_n8136), .b(new_n7299), .O(new_n8137));
  nor2 g07944(.a(new_n8137), .b(new_n8134), .O(new_n8138));
  inv1 g07945(.a(new_n8138), .O(new_n8139));
  nor2 g07946(.a(new_n8139), .b(new_n7980), .O(new_n8140));
  inv1 g07947(.a(new_n7980), .O(new_n8141));
  nor2 g07948(.a(new_n8138), .b(new_n8141), .O(new_n8142));
  nor2 g07949(.a(new_n8142), .b(new_n8140), .O(new_n8143));
  nor2 g07950(.a(new_n6958), .b(new_n214), .O(new_n8144));
  inv1 g07951(.a(new_n8144), .O(new_n8145));
  nor2 g07952(.a(new_n3870), .b(new_n941), .O(new_n8146));
  nor2 g07953(.a(new_n3722), .b(new_n1086), .O(new_n8147));
  nor2 g07954(.a(new_n8147), .b(new_n8146), .O(new_n8148));
  nor2 g07955(.a(new_n3870), .b(new_n1086), .O(new_n8149));
  inv1 g07956(.a(new_n8149), .O(new_n8150));
  nor2 g07957(.a(new_n8150), .b(new_n8023), .O(new_n8151));
  nor2 g07958(.a(new_n8151), .b(new_n8148), .O(new_n8152));
  nor2 g07959(.a(new_n8152), .b(new_n8145), .O(new_n8153));
  inv1 g07960(.a(new_n8152), .O(new_n8154));
  nor2 g07961(.a(new_n8154), .b(new_n8144), .O(new_n8155));
  nor2 g07962(.a(new_n8155), .b(new_n8153), .O(new_n8156));
  nor2 g07963(.a(new_n8156), .b(new_n8143), .O(new_n8157));
  inv1 g07964(.a(new_n8143), .O(new_n8158));
  inv1 g07965(.a(new_n8156), .O(new_n8159));
  nor2 g07966(.a(new_n8159), .b(new_n8158), .O(new_n8160));
  nor2 g07967(.a(new_n8160), .b(new_n8157), .O(new_n8161));
  nor2 g07968(.a(new_n8161), .b(new_n8132), .O(new_n8162));
  inv1 g07969(.a(new_n8161), .O(new_n8163));
  nor2 g07970(.a(new_n8163), .b(new_n8131), .O(new_n8164));
  nor2 g07971(.a(new_n8164), .b(new_n8162), .O(new_n8165));
  nor2 g07972(.a(new_n8165), .b(new_n8119), .O(new_n8166));
  inv1 g07973(.a(new_n8165), .O(new_n8167));
  nor2 g07974(.a(new_n8167), .b(new_n8118), .O(new_n8168));
  nor2 g07975(.a(new_n8168), .b(new_n8166), .O(new_n8169));
  inv1 g07976(.a(\a[53] ), .O(new_n8170));
  nor2 g07977(.a(new_n8170), .b(new_n198), .O(new_n8171));
  inv1 g07978(.a(new_n8171), .O(new_n8172));
  nor2 g07979(.a(new_n6893), .b(new_n229), .O(new_n8173));
  nor2 g07980(.a(new_n4093), .b(new_n847), .O(new_n8174));
  nor2 g07981(.a(new_n8174), .b(new_n8173), .O(new_n8175));
  nor2 g07982(.a(new_n6893), .b(new_n847), .O(new_n8176));
  inv1 g07983(.a(new_n8176), .O(new_n8177));
  nor2 g07984(.a(new_n8177), .b(new_n5161), .O(new_n8178));
  nor2 g07985(.a(new_n8178), .b(new_n8175), .O(new_n8179));
  nor2 g07986(.a(new_n8179), .b(new_n8172), .O(new_n8180));
  inv1 g07987(.a(new_n8179), .O(new_n8181));
  nor2 g07988(.a(new_n8181), .b(new_n8171), .O(new_n8182));
  nor2 g07989(.a(new_n8182), .b(new_n8180), .O(new_n8183));
  nor2 g07990(.a(new_n6570), .b(new_n257), .O(new_n8184));
  inv1 g07991(.a(new_n8184), .O(new_n8185));
  nor2 g07992(.a(new_n4366), .b(new_n800), .O(new_n8186));
  nor2 g07993(.a(new_n6274), .b(new_n295), .O(new_n8187));
  nor2 g07994(.a(new_n8187), .b(new_n8186), .O(new_n8188));
  inv1 g07995(.a(new_n8186), .O(new_n8189));
  inv1 g07996(.a(new_n8187), .O(new_n8190));
  nor2 g07997(.a(new_n8190), .b(new_n8189), .O(new_n8191));
  nor2 g07998(.a(new_n8191), .b(new_n8188), .O(new_n8192));
  nor2 g07999(.a(new_n8192), .b(new_n8185), .O(new_n8193));
  inv1 g08000(.a(new_n8192), .O(new_n8194));
  nor2 g08001(.a(new_n8194), .b(new_n8184), .O(new_n8195));
  nor2 g08002(.a(new_n8195), .b(new_n8193), .O(new_n8196));
  nor2 g08003(.a(new_n5796), .b(new_n363), .O(new_n8197));
  nor2 g08004(.a(new_n4425), .b(new_n699), .O(new_n8198));
  nor2 g08005(.a(new_n8198), .b(new_n8197), .O(new_n8199));
  nor2 g08006(.a(new_n5796), .b(new_n699), .O(new_n8200));
  inv1 g08007(.a(new_n8200), .O(new_n8201));
  nor2 g08008(.a(new_n8201), .b(new_n6677), .O(new_n8202));
  nor2 g08009(.a(new_n8202), .b(new_n8199), .O(new_n8203));
  nor2 g08010(.a(new_n8203), .b(new_n7831), .O(new_n8204));
  inv1 g08011(.a(new_n8203), .O(new_n8205));
  nor2 g08012(.a(new_n8205), .b(new_n7830), .O(new_n8206));
  nor2 g08013(.a(new_n8206), .b(new_n8204), .O(new_n8207));
  nor2 g08014(.a(new_n8207), .b(new_n8196), .O(new_n8208));
  inv1 g08015(.a(new_n8196), .O(new_n8209));
  inv1 g08016(.a(new_n8207), .O(new_n8210));
  nor2 g08017(.a(new_n8210), .b(new_n8209), .O(new_n8211));
  nor2 g08018(.a(new_n8211), .b(new_n8208), .O(new_n8212));
  inv1 g08019(.a(new_n8212), .O(new_n8213));
  nor2 g08020(.a(new_n8213), .b(new_n8183), .O(new_n8214));
  inv1 g08021(.a(new_n8183), .O(new_n8215));
  nor2 g08022(.a(new_n8212), .b(new_n8215), .O(new_n8216));
  nor2 g08023(.a(new_n8216), .b(new_n8214), .O(new_n8217));
  nor2 g08024(.a(new_n8217), .b(new_n8169), .O(new_n8218));
  inv1 g08025(.a(new_n8169), .O(new_n8219));
  inv1 g08026(.a(new_n8217), .O(new_n8220));
  nor2 g08027(.a(new_n8220), .b(new_n8219), .O(new_n8221));
  nor2 g08028(.a(new_n8221), .b(new_n8218), .O(new_n8222));
  inv1 g08029(.a(new_n8222), .O(new_n8223));
  nor2 g08030(.a(new_n7999), .b(new_n7994), .O(new_n8224));
  inv1 g08031(.a(new_n8224), .O(new_n8225));
  nor2 g08032(.a(new_n5178), .b(new_n502), .O(new_n8226));
  inv1 g08033(.a(new_n8226), .O(new_n8227));
  nor2 g08034(.a(new_n2184), .b(new_n2121), .O(new_n8228));
  nor2 g08035(.a(new_n2433), .b(new_n1903), .O(new_n8229));
  nor2 g08036(.a(new_n8229), .b(new_n8228), .O(new_n8230));
  nor2 g08037(.a(new_n2433), .b(new_n2121), .O(new_n8231));
  inv1 g08038(.a(new_n8231), .O(new_n8232));
  nor2 g08039(.a(new_n8232), .b(new_n7615), .O(new_n8233));
  nor2 g08040(.a(new_n8233), .b(new_n8230), .O(new_n8234));
  nor2 g08041(.a(new_n8234), .b(new_n8227), .O(new_n8235));
  inv1 g08042(.a(new_n8234), .O(new_n8236));
  nor2 g08043(.a(new_n8236), .b(new_n8226), .O(new_n8237));
  nor2 g08044(.a(new_n8237), .b(new_n8235), .O(new_n8238));
  inv1 g08045(.a(new_n8238), .O(new_n8239));
  nor2 g08046(.a(new_n4682), .b(new_n613), .O(new_n8240));
  nor2 g08047(.a(new_n5393), .b(new_n438), .O(new_n8241));
  nor2 g08048(.a(new_n8241), .b(new_n7640), .O(new_n8242));
  inv1 g08049(.a(new_n7638), .O(new_n8243));
  nor2 g08050(.a(new_n5393), .b(new_n569), .O(new_n8244));
  inv1 g08051(.a(new_n8244), .O(new_n8245));
  nor2 g08052(.a(new_n8245), .b(new_n8243), .O(new_n8246));
  nor2 g08053(.a(new_n8246), .b(new_n8242), .O(new_n8247));
  inv1 g08054(.a(new_n8247), .O(new_n8248));
  nor2 g08055(.a(new_n8248), .b(new_n8240), .O(new_n8249));
  inv1 g08056(.a(new_n8240), .O(new_n8250));
  nor2 g08057(.a(new_n8247), .b(new_n8250), .O(new_n8251));
  nor2 g08058(.a(new_n8251), .b(new_n8249), .O(new_n8252));
  nor2 g08059(.a(new_n2826), .b(new_n1493), .O(new_n8253));
  inv1 g08060(.a(new_n8253), .O(new_n8254));
  nor2 g08061(.a(new_n2660), .b(new_n1647), .O(new_n8255));
  nor2 g08062(.a(new_n8255), .b(new_n7889), .O(new_n8256));
  nor2 g08063(.a(new_n2660), .b(new_n1736), .O(new_n8257));
  inv1 g08064(.a(new_n8257), .O(new_n8258));
  nor2 g08065(.a(new_n8258), .b(new_n7567), .O(new_n8259));
  nor2 g08066(.a(new_n8259), .b(new_n8256), .O(new_n8260));
  nor2 g08067(.a(new_n8260), .b(new_n8254), .O(new_n8261));
  inv1 g08068(.a(new_n8260), .O(new_n8262));
  nor2 g08069(.a(new_n8262), .b(new_n8253), .O(new_n8263));
  nor2 g08070(.a(new_n8263), .b(new_n8261), .O(new_n8264));
  nor2 g08071(.a(new_n8264), .b(new_n8252), .O(new_n8265));
  inv1 g08072(.a(new_n8252), .O(new_n8266));
  inv1 g08073(.a(new_n8264), .O(new_n8267));
  nor2 g08074(.a(new_n8267), .b(new_n8266), .O(new_n8268));
  nor2 g08075(.a(new_n8268), .b(new_n8265), .O(new_n8269));
  nor2 g08076(.a(new_n8269), .b(new_n8239), .O(new_n8270));
  inv1 g08077(.a(new_n8269), .O(new_n8271));
  nor2 g08078(.a(new_n8271), .b(new_n8238), .O(new_n8272));
  nor2 g08079(.a(new_n8272), .b(new_n8270), .O(new_n8273));
  nor2 g08080(.a(new_n8273), .b(new_n8225), .O(new_n8274));
  inv1 g08081(.a(new_n8273), .O(new_n8275));
  nor2 g08082(.a(new_n8275), .b(new_n8224), .O(new_n8276));
  nor2 g08083(.a(new_n8276), .b(new_n8274), .O(new_n8277));
  inv1 g08084(.a(new_n8277), .O(new_n8278));
  nor2 g08085(.a(new_n8084), .b(new_n8081), .O(new_n8279));
  nor2 g08086(.a(new_n8279), .b(new_n8278), .O(new_n8280));
  inv1 g08087(.a(new_n8279), .O(new_n8281));
  nor2 g08088(.a(new_n8281), .b(new_n8277), .O(new_n8282));
  nor2 g08089(.a(new_n8282), .b(new_n8280), .O(new_n8283));
  inv1 g08090(.a(new_n8283), .O(new_n8284));
  nor2 g08091(.a(new_n8284), .b(new_n8223), .O(new_n8285));
  nor2 g08092(.a(new_n8283), .b(new_n8222), .O(new_n8286));
  nor2 g08093(.a(new_n8286), .b(new_n8285), .O(new_n8287));
  inv1 g08094(.a(new_n8287), .O(new_n8288));
  nor2 g08095(.a(new_n8288), .b(new_n8117), .O(new_n8289));
  inv1 g08096(.a(new_n8117), .O(new_n8290));
  nor2 g08097(.a(new_n8287), .b(new_n8290), .O(new_n8291));
  nor2 g08098(.a(new_n8291), .b(new_n8289), .O(new_n8292));
  inv1 g08099(.a(new_n8292), .O(new_n8293));
  nor2 g08100(.a(new_n8293), .b(new_n8116), .O(new_n8294));
  inv1 g08101(.a(new_n8116), .O(new_n8295));
  nor2 g08102(.a(new_n8292), .b(new_n8295), .O(new_n8296));
  nor2 g08103(.a(new_n8296), .b(new_n8294), .O(new_n8297));
  inv1 g08104(.a(new_n8297), .O(new_n8298));
  nor2 g08105(.a(new_n8004), .b(new_n7972), .O(new_n8299));
  inv1 g08106(.a(new_n8299), .O(new_n8300));
  nor2 g08107(.a(new_n7957), .b(new_n7950), .O(new_n8301));
  nor2 g08108(.a(new_n8031), .b(new_n8022), .O(new_n8302));
  nor2 g08109(.a(new_n8302), .b(new_n8301), .O(new_n8303));
  inv1 g08110(.a(new_n8301), .O(new_n8304));
  inv1 g08111(.a(new_n8302), .O(new_n8305));
  nor2 g08112(.a(new_n8305), .b(new_n8304), .O(new_n8306));
  nor2 g08113(.a(new_n8306), .b(new_n8303), .O(new_n8307));
  nor2 g08114(.a(new_n7895), .b(new_n7887), .O(new_n8308));
  nor2 g08115(.a(new_n8308), .b(new_n8307), .O(new_n8309));
  inv1 g08116(.a(new_n8307), .O(new_n8310));
  inv1 g08117(.a(new_n8308), .O(new_n8311));
  nor2 g08118(.a(new_n8311), .b(new_n8310), .O(new_n8312));
  nor2 g08119(.a(new_n8312), .b(new_n8309), .O(new_n8313));
  inv1 g08120(.a(new_n8313), .O(new_n8314));
  nor2 g08121(.a(new_n7912), .b(new_n7897), .O(new_n8315));
  inv1 g08122(.a(new_n8315), .O(new_n8316));
  nor2 g08123(.a(new_n8036), .b(new_n8019), .O(new_n8317));
  inv1 g08124(.a(new_n8317), .O(new_n8318));
  nor2 g08125(.a(new_n8318), .b(new_n8316), .O(new_n8319));
  nor2 g08126(.a(new_n8317), .b(new_n8315), .O(new_n8320));
  nor2 g08127(.a(new_n8320), .b(new_n8319), .O(new_n8321));
  inv1 g08128(.a(new_n8321), .O(new_n8322));
  nor2 g08129(.a(new_n8322), .b(new_n8314), .O(new_n8323));
  nor2 g08130(.a(new_n8321), .b(new_n8313), .O(new_n8324));
  nor2 g08131(.a(new_n8324), .b(new_n8323), .O(new_n8325));
  inv1 g08132(.a(new_n8325), .O(new_n8326));
  nor2 g08133(.a(new_n7859), .b(new_n7852), .O(new_n8327));
  nor2 g08134(.a(new_n7880), .b(new_n7873), .O(new_n8328));
  nor2 g08135(.a(new_n8328), .b(new_n8327), .O(new_n8329));
  inv1 g08136(.a(new_n8327), .O(new_n8330));
  inv1 g08137(.a(new_n8328), .O(new_n8331));
  nor2 g08138(.a(new_n8331), .b(new_n8330), .O(new_n8332));
  nor2 g08139(.a(new_n8332), .b(new_n8329), .O(new_n8333));
  nor2 g08140(.a(new_n7836), .b(new_n7829), .O(new_n8334));
  nor2 g08141(.a(new_n8334), .b(new_n8333), .O(new_n8335));
  inv1 g08142(.a(new_n8333), .O(new_n8336));
  inv1 g08143(.a(new_n8334), .O(new_n8337));
  nor2 g08144(.a(new_n8337), .b(new_n8336), .O(new_n8338));
  nor2 g08145(.a(new_n8338), .b(new_n8335), .O(new_n8339));
  inv1 g08146(.a(new_n8339), .O(new_n8340));
  nor2 g08147(.a(new_n7867), .b(new_n7861), .O(new_n8341));
  nor2 g08148(.a(new_n2367), .b(new_n8026), .O(new_n8342));
  nor2 g08149(.a(new_n8026), .b(new_n194), .O(new_n8343));
  nor2 g08150(.a(new_n8343), .b(\a[27] ), .O(new_n8344));
  nor2 g08151(.a(new_n8344), .b(new_n8342), .O(new_n8345));
  nor2 g08152(.a(new_n7846), .b(new_n7841), .O(new_n8346));
  nor2 g08153(.a(new_n8346), .b(new_n8345), .O(new_n8347));
  inv1 g08154(.a(new_n8345), .O(new_n8348));
  inv1 g08155(.a(new_n8346), .O(new_n8349));
  nor2 g08156(.a(new_n8349), .b(new_n8348), .O(new_n8350));
  nor2 g08157(.a(new_n8350), .b(new_n8347), .O(new_n8351));
  inv1 g08158(.a(new_n8351), .O(new_n8352));
  nor2 g08159(.a(new_n7910), .b(new_n7905), .O(new_n8353));
  inv1 g08160(.a(new_n8353), .O(new_n8354));
  nor2 g08161(.a(new_n8354), .b(new_n8352), .O(new_n8355));
  nor2 g08162(.a(new_n8353), .b(new_n8351), .O(new_n8356));
  nor2 g08163(.a(new_n8356), .b(new_n8355), .O(new_n8357));
  inv1 g08164(.a(new_n8357), .O(new_n8358));
  nor2 g08165(.a(new_n8358), .b(new_n8341), .O(new_n8359));
  inv1 g08166(.a(new_n8341), .O(new_n8360));
  nor2 g08167(.a(new_n8357), .b(new_n8360), .O(new_n8361));
  nor2 g08168(.a(new_n8361), .b(new_n8359), .O(new_n8362));
  inv1 g08169(.a(new_n8362), .O(new_n8363));
  nor2 g08170(.a(new_n8363), .b(new_n8340), .O(new_n8364));
  nor2 g08171(.a(new_n8362), .b(new_n8339), .O(new_n8365));
  nor2 g08172(.a(new_n8365), .b(new_n8364), .O(new_n8366));
  inv1 g08173(.a(new_n8366), .O(new_n8367));
  nor2 g08174(.a(new_n8367), .b(new_n8326), .O(new_n8368));
  nor2 g08175(.a(new_n8366), .b(new_n8325), .O(new_n8369));
  nor2 g08176(.a(new_n8369), .b(new_n8368), .O(new_n8370));
  nor2 g08177(.a(new_n8370), .b(new_n8300), .O(new_n8371));
  inv1 g08178(.a(new_n8370), .O(new_n8372));
  nor2 g08179(.a(new_n8372), .b(new_n8299), .O(new_n8373));
  nor2 g08180(.a(new_n8373), .b(new_n8371), .O(new_n8374));
  inv1 g08181(.a(new_n8374), .O(new_n8375));
  nor2 g08182(.a(new_n7922), .b(new_n7919), .O(new_n8376));
  nor2 g08183(.a(new_n8061), .b(new_n8055), .O(new_n8377));
  inv1 g08184(.a(new_n8377), .O(new_n8378));
  nor2 g08185(.a(new_n7989), .b(new_n7983), .O(new_n8379));
  inv1 g08186(.a(new_n8379), .O(new_n8380));
  nor2 g08187(.a(new_n8380), .b(new_n8378), .O(new_n8381));
  nor2 g08188(.a(new_n8379), .b(new_n8377), .O(new_n8382));
  nor2 g08189(.a(new_n8382), .b(new_n8381), .O(new_n8383));
  nor2 g08190(.a(new_n8075), .b(new_n8069), .O(new_n8384));
  inv1 g08191(.a(new_n8384), .O(new_n8385));
  nor2 g08192(.a(new_n8385), .b(new_n8383), .O(new_n8386));
  inv1 g08193(.a(new_n8383), .O(new_n8387));
  nor2 g08194(.a(new_n8384), .b(new_n8387), .O(new_n8388));
  nor2 g08195(.a(new_n8388), .b(new_n8386), .O(new_n8389));
  nor2 g08196(.a(new_n8046), .b(new_n8040), .O(new_n8390));
  inv1 g08197(.a(new_n8390), .O(new_n8391));
  nor2 g08198(.a(new_n8391), .b(new_n8389), .O(new_n8392));
  inv1 g08199(.a(new_n8389), .O(new_n8393));
  nor2 g08200(.a(new_n8390), .b(new_n8393), .O(new_n8394));
  nor2 g08201(.a(new_n8394), .b(new_n8392), .O(new_n8395));
  inv1 g08202(.a(new_n8395), .O(new_n8396));
  nor2 g08203(.a(new_n8396), .b(new_n8376), .O(new_n8397));
  inv1 g08204(.a(new_n8376), .O(new_n8398));
  nor2 g08205(.a(new_n8395), .b(new_n8398), .O(new_n8399));
  nor2 g08206(.a(new_n8399), .b(new_n8397), .O(new_n8400));
  nor2 g08207(.a(new_n7933), .b(new_n7927), .O(new_n8401));
  inv1 g08208(.a(new_n8401), .O(new_n8402));
  nor2 g08209(.a(new_n8402), .b(new_n8400), .O(new_n8403));
  inv1 g08210(.a(new_n8400), .O(new_n8404));
  nor2 g08211(.a(new_n8401), .b(new_n8404), .O(new_n8405));
  nor2 g08212(.a(new_n8405), .b(new_n8403), .O(new_n8406));
  inv1 g08213(.a(new_n8406), .O(new_n8407));
  nor2 g08214(.a(new_n8407), .b(new_n8375), .O(new_n8408));
  nor2 g08215(.a(new_n8406), .b(new_n8374), .O(new_n8409));
  nor2 g08216(.a(new_n8409), .b(new_n8408), .O(new_n8410));
  inv1 g08217(.a(new_n8410), .O(new_n8411));
  nor2 g08218(.a(new_n8411), .b(new_n8298), .O(new_n8412));
  nor2 g08219(.a(new_n8410), .b(new_n8297), .O(new_n8413));
  nor2 g08220(.a(new_n8413), .b(new_n8412), .O(new_n8414));
  inv1 g08221(.a(new_n8414), .O(new_n8415));
  nor2 g08222(.a(new_n8415), .b(new_n8115), .O(new_n8416));
  inv1 g08223(.a(new_n8115), .O(new_n8417));
  nor2 g08224(.a(new_n8414), .b(new_n8417), .O(new_n8418));
  nor2 g08225(.a(new_n8418), .b(new_n8416), .O(new_n8419));
  inv1 g08226(.a(new_n8419), .O(new_n8420));
  nor2 g08227(.a(new_n8112), .b(new_n8104), .O(new_n8421));
  nor2 g08228(.a(new_n8421), .b(new_n8420), .O(new_n8422));
  inv1 g08229(.a(new_n8421), .O(new_n8423));
  nor2 g08230(.a(new_n8423), .b(new_n8419), .O(new_n8424));
  nor2 g08231(.a(new_n8424), .b(new_n8422), .O(new_n8425));
  inv1 g08232(.a(new_n8425), .O(\asquared[54] ));
  nor2 g08233(.a(new_n8412), .b(new_n8294), .O(new_n8427));
  nor2 g08234(.a(new_n8408), .b(new_n8405), .O(new_n8428));
  nor2 g08235(.a(new_n8373), .b(new_n8368), .O(new_n8429));
  inv1 g08236(.a(new_n8429), .O(new_n8430));
  nor2 g08237(.a(new_n8397), .b(new_n8394), .O(new_n8431));
  inv1 g08238(.a(new_n8431), .O(new_n8432));
  nor2 g08239(.a(new_n8432), .b(new_n8430), .O(new_n8433));
  nor2 g08240(.a(new_n8431), .b(new_n8429), .O(new_n8434));
  nor2 g08241(.a(new_n8434), .b(new_n8433), .O(new_n8435));
  inv1 g08242(.a(new_n8435), .O(new_n8436));
  nor2 g08243(.a(new_n8364), .b(new_n8359), .O(new_n8437));
  nor2 g08244(.a(new_n8323), .b(new_n8320), .O(new_n8438));
  nor2 g08245(.a(new_n3722), .b(new_n1199), .O(new_n8439));
  nor2 g08246(.a(new_n3057), .b(new_n1493), .O(new_n8440));
  nor2 g08247(.a(new_n8440), .b(new_n8124), .O(new_n8441));
  nor2 g08248(.a(new_n3231), .b(new_n1493), .O(new_n8442));
  inv1 g08249(.a(new_n8442), .O(new_n8443));
  nor2 g08250(.a(new_n8443), .b(new_n7876), .O(new_n8444));
  nor2 g08251(.a(new_n8444), .b(new_n8441), .O(new_n8445));
  inv1 g08252(.a(new_n8445), .O(new_n8446));
  nor2 g08253(.a(new_n8446), .b(new_n8439), .O(new_n8447));
  inv1 g08254(.a(new_n8439), .O(new_n8448));
  nor2 g08255(.a(new_n8445), .b(new_n8448), .O(new_n8449));
  nor2 g08256(.a(new_n8449), .b(new_n8447), .O(new_n8450));
  nor2 g08257(.a(new_n2826), .b(new_n1647), .O(new_n8451));
  inv1 g08258(.a(new_n8451), .O(new_n8452));
  nor2 g08259(.a(new_n2506), .b(new_n1903), .O(new_n8453));
  nor2 g08260(.a(new_n8453), .b(new_n8257), .O(new_n8454));
  nor2 g08261(.a(new_n2660), .b(new_n1903), .O(new_n8455));
  inv1 g08262(.a(new_n8455), .O(new_n8456));
  nor2 g08263(.a(new_n8456), .b(new_n7890), .O(new_n8457));
  nor2 g08264(.a(new_n8457), .b(new_n8454), .O(new_n8458));
  nor2 g08265(.a(new_n8458), .b(new_n8452), .O(new_n8459));
  inv1 g08266(.a(new_n8458), .O(new_n8460));
  nor2 g08267(.a(new_n8460), .b(new_n8451), .O(new_n8461));
  nor2 g08268(.a(new_n8461), .b(new_n8459), .O(new_n8462));
  nor2 g08269(.a(new_n8462), .b(new_n8450), .O(new_n8463));
  inv1 g08270(.a(new_n8450), .O(new_n8464));
  inv1 g08271(.a(new_n8462), .O(new_n8465));
  nor2 g08272(.a(new_n8465), .b(new_n8464), .O(new_n8466));
  nor2 g08273(.a(new_n8466), .b(new_n8463), .O(new_n8467));
  inv1 g08274(.a(new_n8467), .O(new_n8468));
  nor2 g08275(.a(new_n8170), .b(new_n194), .O(new_n8469));
  nor2 g08276(.a(new_n8469), .b(new_n8231), .O(new_n8470));
  inv1 g08277(.a(new_n8469), .O(new_n8471));
  nor2 g08278(.a(new_n8471), .b(new_n8232), .O(new_n8472));
  nor2 g08279(.a(new_n8472), .b(new_n8470), .O(new_n8473));
  inv1 g08280(.a(new_n8473), .O(new_n8474));
  inv1 g08281(.a(new_n8342), .O(new_n8475));
  inv1 g08282(.a(\a[54] ), .O(new_n8476));
  nor2 g08283(.a(new_n8476), .b(new_n198), .O(new_n8477));
  inv1 g08284(.a(new_n8477), .O(new_n8478));
  nor2 g08285(.a(new_n8478), .b(new_n8475), .O(new_n8479));
  nor2 g08286(.a(new_n8477), .b(new_n8342), .O(new_n8480));
  nor2 g08287(.a(new_n8480), .b(new_n8479), .O(new_n8481));
  inv1 g08288(.a(new_n8481), .O(new_n8482));
  nor2 g08289(.a(new_n8482), .b(new_n8474), .O(new_n8483));
  nor2 g08290(.a(new_n8481), .b(new_n8473), .O(new_n8484));
  nor2 g08291(.a(new_n8484), .b(new_n8483), .O(new_n8485));
  inv1 g08292(.a(new_n8485), .O(new_n8486));
  nor2 g08293(.a(new_n8486), .b(new_n8468), .O(new_n8487));
  nor2 g08294(.a(new_n8485), .b(new_n8467), .O(new_n8488));
  nor2 g08295(.a(new_n8488), .b(new_n8487), .O(new_n8489));
  inv1 g08296(.a(new_n8489), .O(new_n8490));
  nor2 g08297(.a(new_n8490), .b(new_n8438), .O(new_n8491));
  inv1 g08298(.a(new_n8438), .O(new_n8492));
  nor2 g08299(.a(new_n8489), .b(new_n8492), .O(new_n8493));
  nor2 g08300(.a(new_n8493), .b(new_n8491), .O(new_n8494));
  inv1 g08301(.a(new_n8494), .O(new_n8495));
  nor2 g08302(.a(new_n8495), .b(new_n8437), .O(new_n8496));
  inv1 g08303(.a(new_n8437), .O(new_n8497));
  nor2 g08304(.a(new_n8494), .b(new_n8497), .O(new_n8498));
  nor2 g08305(.a(new_n8498), .b(new_n8496), .O(new_n8499));
  inv1 g08306(.a(new_n8499), .O(new_n8500));
  nor2 g08307(.a(new_n8500), .b(new_n8436), .O(new_n8501));
  nor2 g08308(.a(new_n8499), .b(new_n8435), .O(new_n8502));
  nor2 g08309(.a(new_n8502), .b(new_n8501), .O(new_n8503));
  inv1 g08310(.a(new_n8503), .O(new_n8504));
  nor2 g08311(.a(new_n8504), .b(new_n8428), .O(new_n8505));
  inv1 g08312(.a(new_n8428), .O(new_n8506));
  nor2 g08313(.a(new_n8503), .b(new_n8506), .O(new_n8507));
  nor2 g08314(.a(new_n8507), .b(new_n8505), .O(new_n8508));
  inv1 g08315(.a(new_n8508), .O(new_n8509));
  nor2 g08316(.a(new_n8289), .b(new_n8285), .O(new_n8510));
  inv1 g08317(.a(new_n8510), .O(new_n8511));
  nor2 g08318(.a(new_n8338), .b(new_n8332), .O(new_n8512));
  inv1 g08319(.a(new_n8512), .O(new_n8513));
  nor2 g08320(.a(new_n8312), .b(new_n8306), .O(new_n8514));
  inv1 g08321(.a(new_n8514), .O(new_n8515));
  nor2 g08322(.a(new_n8515), .b(new_n8513), .O(new_n8516));
  nor2 g08323(.a(new_n8514), .b(new_n8512), .O(new_n8517));
  nor2 g08324(.a(new_n8517), .b(new_n8516), .O(new_n8518));
  nor2 g08325(.a(new_n8355), .b(new_n8350), .O(new_n8519));
  inv1 g08326(.a(new_n8519), .O(new_n8520));
  nor2 g08327(.a(new_n8520), .b(new_n8518), .O(new_n8521));
  inv1 g08328(.a(new_n8518), .O(new_n8522));
  nor2 g08329(.a(new_n8519), .b(new_n8522), .O(new_n8523));
  nor2 g08330(.a(new_n8523), .b(new_n8521), .O(new_n8524));
  inv1 g08331(.a(new_n8524), .O(new_n8525));
  nor2 g08332(.a(new_n8221), .b(new_n8168), .O(new_n8526));
  nor2 g08333(.a(new_n8526), .b(new_n8525), .O(new_n8527));
  inv1 g08334(.a(new_n8526), .O(new_n8528));
  nor2 g08335(.a(new_n8528), .b(new_n8524), .O(new_n8529));
  nor2 g08336(.a(new_n8529), .b(new_n8527), .O(new_n8530));
  inv1 g08337(.a(new_n8530), .O(new_n8531));
  nor2 g08338(.a(new_n8195), .b(new_n8188), .O(new_n8532));
  nor2 g08339(.a(new_n8182), .b(new_n8175), .O(new_n8533));
  nor2 g08340(.a(new_n8533), .b(new_n8532), .O(new_n8534));
  inv1 g08341(.a(new_n8532), .O(new_n8535));
  inv1 g08342(.a(new_n8533), .O(new_n8536));
  nor2 g08343(.a(new_n8536), .b(new_n8535), .O(new_n8537));
  nor2 g08344(.a(new_n8537), .b(new_n8534), .O(new_n8538));
  nor2 g08345(.a(new_n8237), .b(new_n8230), .O(new_n8539));
  nor2 g08346(.a(new_n8539), .b(new_n8538), .O(new_n8540));
  inv1 g08347(.a(new_n8538), .O(new_n8541));
  inv1 g08348(.a(new_n8539), .O(new_n8542));
  nor2 g08349(.a(new_n8542), .b(new_n8541), .O(new_n8543));
  nor2 g08350(.a(new_n8543), .b(new_n8540), .O(new_n8544));
  inv1 g08351(.a(new_n8544), .O(new_n8545));
  nor2 g08352(.a(new_n8155), .b(new_n8148), .O(new_n8546));
  nor2 g08353(.a(new_n8130), .b(new_n8123), .O(new_n8547));
  nor2 g08354(.a(new_n8547), .b(new_n8546), .O(new_n8548));
  inv1 g08355(.a(new_n8546), .O(new_n8549));
  inv1 g08356(.a(new_n8547), .O(new_n8550));
  nor2 g08357(.a(new_n8550), .b(new_n8549), .O(new_n8551));
  nor2 g08358(.a(new_n8551), .b(new_n8548), .O(new_n8552));
  nor2 g08359(.a(new_n8263), .b(new_n8256), .O(new_n8553));
  nor2 g08360(.a(new_n8553), .b(new_n8552), .O(new_n8554));
  inv1 g08361(.a(new_n8552), .O(new_n8555));
  inv1 g08362(.a(new_n8553), .O(new_n8556));
  nor2 g08363(.a(new_n8556), .b(new_n8555), .O(new_n8557));
  nor2 g08364(.a(new_n8557), .b(new_n8554), .O(new_n8558));
  nor2 g08365(.a(new_n8214), .b(new_n8208), .O(new_n8559));
  inv1 g08366(.a(new_n8559), .O(new_n8560));
  nor2 g08367(.a(new_n8560), .b(new_n8558), .O(new_n8561));
  inv1 g08368(.a(new_n8558), .O(new_n8562));
  nor2 g08369(.a(new_n8559), .b(new_n8562), .O(new_n8563));
  nor2 g08370(.a(new_n8563), .b(new_n8561), .O(new_n8564));
  inv1 g08371(.a(new_n8564), .O(new_n8565));
  nor2 g08372(.a(new_n8565), .b(new_n8545), .O(new_n8566));
  nor2 g08373(.a(new_n8564), .b(new_n8544), .O(new_n8567));
  nor2 g08374(.a(new_n8567), .b(new_n8566), .O(new_n8568));
  inv1 g08375(.a(new_n8568), .O(new_n8569));
  nor2 g08376(.a(new_n8569), .b(new_n8531), .O(new_n8570));
  nor2 g08377(.a(new_n8568), .b(new_n8530), .O(new_n8571));
  nor2 g08378(.a(new_n8571), .b(new_n8570), .O(new_n8572));
  nor2 g08379(.a(new_n8572), .b(new_n8511), .O(new_n8573));
  inv1 g08380(.a(new_n8572), .O(new_n8574));
  nor2 g08381(.a(new_n8574), .b(new_n8510), .O(new_n8575));
  nor2 g08382(.a(new_n8575), .b(new_n8573), .O(new_n8576));
  inv1 g08383(.a(new_n8576), .O(new_n8577));
  nor2 g08384(.a(new_n8388), .b(new_n8382), .O(new_n8578));
  inv1 g08385(.a(new_n8578), .O(new_n8579));
  nor2 g08386(.a(new_n4093), .b(new_n941), .O(new_n8580));
  inv1 g08387(.a(new_n8580), .O(new_n8581));
  nor2 g08388(.a(new_n6893), .b(new_n257), .O(new_n8582));
  nor2 g08389(.a(new_n4366), .b(new_n847), .O(new_n8583));
  nor2 g08390(.a(new_n8583), .b(new_n8582), .O(new_n8584));
  nor2 g08391(.a(new_n8177), .b(new_n5662), .O(new_n8585));
  nor2 g08392(.a(new_n8585), .b(new_n8584), .O(new_n8586));
  nor2 g08393(.a(new_n8586), .b(new_n8581), .O(new_n8587));
  inv1 g08394(.a(new_n8586), .O(new_n8588));
  nor2 g08395(.a(new_n8588), .b(new_n8580), .O(new_n8589));
  nor2 g08396(.a(new_n8589), .b(new_n8587), .O(new_n8590));
  inv1 g08397(.a(new_n8590), .O(new_n8591));
  nor2 g08398(.a(new_n5178), .b(new_n569), .O(new_n8592));
  nor2 g08399(.a(new_n5393), .b(new_n502), .O(new_n8593));
  nor2 g08400(.a(new_n8593), .b(new_n8592), .O(new_n8594));
  nor2 g08401(.a(new_n8245), .b(new_n8227), .O(new_n8595));
  nor2 g08402(.a(new_n8595), .b(new_n8594), .O(new_n8596));
  nor2 g08403(.a(new_n8596), .b(new_n7334), .O(new_n8597));
  inv1 g08404(.a(new_n8596), .O(new_n8598));
  nor2 g08405(.a(new_n8598), .b(new_n7333), .O(new_n8599));
  nor2 g08406(.a(new_n8599), .b(new_n8597), .O(new_n8600));
  nor2 g08407(.a(new_n3533), .b(new_n1297), .O(new_n8601));
  inv1 g08408(.a(new_n8601), .O(new_n8602));
  nor2 g08409(.a(new_n6958), .b(new_n229), .O(new_n8603));
  nor2 g08410(.a(new_n8603), .b(new_n8149), .O(new_n8604));
  inv1 g08411(.a(new_n8603), .O(new_n8605));
  nor2 g08412(.a(new_n8605), .b(new_n8150), .O(new_n8606));
  nor2 g08413(.a(new_n8606), .b(new_n8604), .O(new_n8607));
  nor2 g08414(.a(new_n8607), .b(new_n8602), .O(new_n8608));
  inv1 g08415(.a(new_n8607), .O(new_n8609));
  nor2 g08416(.a(new_n8609), .b(new_n8601), .O(new_n8610));
  nor2 g08417(.a(new_n8610), .b(new_n8608), .O(new_n8611));
  nor2 g08418(.a(new_n8611), .b(new_n8600), .O(new_n8612));
  inv1 g08419(.a(new_n8600), .O(new_n8613));
  inv1 g08420(.a(new_n8611), .O(new_n8614));
  nor2 g08421(.a(new_n8614), .b(new_n8613), .O(new_n8615));
  nor2 g08422(.a(new_n8615), .b(new_n8612), .O(new_n8616));
  nor2 g08423(.a(new_n8616), .b(new_n8591), .O(new_n8617));
  inv1 g08424(.a(new_n8616), .O(new_n8618));
  nor2 g08425(.a(new_n8618), .b(new_n8590), .O(new_n8619));
  nor2 g08426(.a(new_n8619), .b(new_n8617), .O(new_n8620));
  nor2 g08427(.a(new_n8620), .b(new_n8579), .O(new_n8621));
  inv1 g08428(.a(new_n8620), .O(new_n8622));
  nor2 g08429(.a(new_n8622), .b(new_n8578), .O(new_n8623));
  nor2 g08430(.a(new_n8623), .b(new_n8621), .O(new_n8624));
  nor2 g08431(.a(new_n8026), .b(new_n196), .O(new_n8625));
  nor2 g08432(.a(new_n7294), .b(new_n214), .O(new_n8626));
  nor2 g08433(.a(new_n8626), .b(new_n8135), .O(new_n8627));
  nor2 g08434(.a(new_n7537), .b(new_n214), .O(new_n8628));
  inv1 g08435(.a(new_n8628), .O(new_n8629));
  nor2 g08436(.a(new_n8629), .b(new_n7952), .O(new_n8630));
  nor2 g08437(.a(new_n8630), .b(new_n8627), .O(new_n8631));
  inv1 g08438(.a(new_n8631), .O(new_n8632));
  nor2 g08439(.a(new_n8632), .b(new_n8625), .O(new_n8633));
  inv1 g08440(.a(new_n8625), .O(new_n8634));
  nor2 g08441(.a(new_n8631), .b(new_n8634), .O(new_n8635));
  nor2 g08442(.a(new_n8635), .b(new_n8633), .O(new_n8636));
  nor2 g08443(.a(new_n6570), .b(new_n295), .O(new_n8637));
  inv1 g08444(.a(new_n8637), .O(new_n8638));
  nor2 g08445(.a(new_n4425), .b(new_n800), .O(new_n8639));
  nor2 g08446(.a(new_n6274), .b(new_n322), .O(new_n8640));
  nor2 g08447(.a(new_n8640), .b(new_n8639), .O(new_n8641));
  inv1 g08448(.a(new_n8639), .O(new_n8642));
  inv1 g08449(.a(new_n8640), .O(new_n8643));
  nor2 g08450(.a(new_n8643), .b(new_n8642), .O(new_n8644));
  nor2 g08451(.a(new_n8644), .b(new_n8641), .O(new_n8645));
  nor2 g08452(.a(new_n8645), .b(new_n8638), .O(new_n8646));
  inv1 g08453(.a(new_n8645), .O(new_n8647));
  nor2 g08454(.a(new_n8647), .b(new_n8637), .O(new_n8648));
  nor2 g08455(.a(new_n8648), .b(new_n8646), .O(new_n8649));
  nor2 g08456(.a(new_n8649), .b(new_n8636), .O(new_n8650));
  inv1 g08457(.a(new_n8636), .O(new_n8651));
  inv1 g08458(.a(new_n8649), .O(new_n8652));
  nor2 g08459(.a(new_n8652), .b(new_n8651), .O(new_n8653));
  nor2 g08460(.a(new_n8653), .b(new_n8650), .O(new_n8654));
  inv1 g08461(.a(new_n8654), .O(new_n8655));
  nor2 g08462(.a(new_n5971), .b(new_n363), .O(new_n8656));
  inv1 g08463(.a(new_n8656), .O(new_n8657));
  nor2 g08464(.a(new_n4682), .b(new_n699), .O(new_n8658));
  nor2 g08465(.a(new_n5796), .b(new_n438), .O(new_n8659));
  nor2 g08466(.a(new_n8659), .b(new_n8658), .O(new_n8660));
  inv1 g08467(.a(new_n7318), .O(new_n8661));
  nor2 g08468(.a(new_n8201), .b(new_n8661), .O(new_n8662));
  nor2 g08469(.a(new_n8662), .b(new_n8660), .O(new_n8663));
  nor2 g08470(.a(new_n8663), .b(new_n8657), .O(new_n8664));
  inv1 g08471(.a(new_n8663), .O(new_n8665));
  nor2 g08472(.a(new_n8665), .b(new_n8656), .O(new_n8666));
  nor2 g08473(.a(new_n8666), .b(new_n8664), .O(new_n8667));
  nor2 g08474(.a(new_n8667), .b(new_n8655), .O(new_n8668));
  inv1 g08475(.a(new_n8667), .O(new_n8669));
  nor2 g08476(.a(new_n8669), .b(new_n8654), .O(new_n8670));
  nor2 g08477(.a(new_n8670), .b(new_n8668), .O(new_n8671));
  nor2 g08478(.a(new_n8671), .b(new_n8624), .O(new_n8672));
  inv1 g08479(.a(new_n8624), .O(new_n8673));
  inv1 g08480(.a(new_n8671), .O(new_n8674));
  nor2 g08481(.a(new_n8674), .b(new_n8673), .O(new_n8675));
  nor2 g08482(.a(new_n8675), .b(new_n8672), .O(new_n8676));
  inv1 g08483(.a(new_n8676), .O(new_n8677));
  nor2 g08484(.a(new_n8280), .b(new_n8276), .O(new_n8678));
  nor2 g08485(.a(new_n8206), .b(new_n8199), .O(new_n8679));
  nor2 g08486(.a(new_n8140), .b(new_n8134), .O(new_n8680));
  nor2 g08487(.a(new_n8680), .b(new_n8679), .O(new_n8681));
  inv1 g08488(.a(new_n8679), .O(new_n8682));
  inv1 g08489(.a(new_n8680), .O(new_n8683));
  nor2 g08490(.a(new_n8683), .b(new_n8682), .O(new_n8684));
  nor2 g08491(.a(new_n8684), .b(new_n8681), .O(new_n8685));
  nor2 g08492(.a(new_n8249), .b(new_n8242), .O(new_n8686));
  nor2 g08493(.a(new_n8686), .b(new_n8685), .O(new_n8687));
  inv1 g08494(.a(new_n8685), .O(new_n8688));
  inv1 g08495(.a(new_n8686), .O(new_n8689));
  nor2 g08496(.a(new_n8689), .b(new_n8688), .O(new_n8690));
  nor2 g08497(.a(new_n8690), .b(new_n8687), .O(new_n8691));
  inv1 g08498(.a(new_n8691), .O(new_n8692));
  nor2 g08499(.a(new_n8272), .b(new_n8265), .O(new_n8693));
  inv1 g08500(.a(new_n8693), .O(new_n8694));
  nor2 g08501(.a(new_n8164), .b(new_n8157), .O(new_n8695));
  inv1 g08502(.a(new_n8695), .O(new_n8696));
  nor2 g08503(.a(new_n8696), .b(new_n8694), .O(new_n8697));
  nor2 g08504(.a(new_n8695), .b(new_n8693), .O(new_n8698));
  nor2 g08505(.a(new_n8698), .b(new_n8697), .O(new_n8699));
  inv1 g08506(.a(new_n8699), .O(new_n8700));
  nor2 g08507(.a(new_n8700), .b(new_n8692), .O(new_n8701));
  nor2 g08508(.a(new_n8699), .b(new_n8691), .O(new_n8702));
  nor2 g08509(.a(new_n8702), .b(new_n8701), .O(new_n8703));
  inv1 g08510(.a(new_n8703), .O(new_n8704));
  nor2 g08511(.a(new_n8704), .b(new_n8678), .O(new_n8705));
  inv1 g08512(.a(new_n8678), .O(new_n8706));
  nor2 g08513(.a(new_n8703), .b(new_n8706), .O(new_n8707));
  nor2 g08514(.a(new_n8707), .b(new_n8705), .O(new_n8708));
  inv1 g08515(.a(new_n8708), .O(new_n8709));
  nor2 g08516(.a(new_n8709), .b(new_n8677), .O(new_n8710));
  nor2 g08517(.a(new_n8708), .b(new_n8676), .O(new_n8711));
  nor2 g08518(.a(new_n8711), .b(new_n8710), .O(new_n8712));
  inv1 g08519(.a(new_n8712), .O(new_n8713));
  nor2 g08520(.a(new_n8713), .b(new_n8577), .O(new_n8714));
  nor2 g08521(.a(new_n8712), .b(new_n8576), .O(new_n8715));
  nor2 g08522(.a(new_n8715), .b(new_n8714), .O(new_n8716));
  inv1 g08523(.a(new_n8716), .O(new_n8717));
  nor2 g08524(.a(new_n8717), .b(new_n8509), .O(new_n8718));
  nor2 g08525(.a(new_n8716), .b(new_n8508), .O(new_n8719));
  nor2 g08526(.a(new_n8719), .b(new_n8718), .O(new_n8720));
  inv1 g08527(.a(new_n8720), .O(new_n8721));
  nor2 g08528(.a(new_n8721), .b(new_n8427), .O(new_n8722));
  inv1 g08529(.a(new_n8427), .O(new_n8723));
  nor2 g08530(.a(new_n8720), .b(new_n8723), .O(new_n8724));
  nor2 g08531(.a(new_n8724), .b(new_n8722), .O(new_n8725));
  nor2 g08532(.a(new_n8422), .b(new_n8418), .O(new_n8726));
  inv1 g08533(.a(new_n8726), .O(new_n8727));
  nor2 g08534(.a(new_n8727), .b(new_n8725), .O(new_n8728));
  inv1 g08535(.a(new_n8725), .O(new_n8729));
  nor2 g08536(.a(new_n8726), .b(new_n8729), .O(new_n8730));
  nor2 g08537(.a(new_n8730), .b(new_n8728), .O(new_n8731));
  inv1 g08538(.a(new_n8731), .O(\asquared[55] ));
  nor2 g08539(.a(new_n8718), .b(new_n8505), .O(new_n8733));
  nor2 g08540(.a(new_n8501), .b(new_n8434), .O(new_n8734));
  inv1 g08541(.a(new_n8734), .O(new_n8735));
  nor2 g08542(.a(new_n8675), .b(new_n8623), .O(new_n8736));
  nor2 g08543(.a(new_n8543), .b(new_n8537), .O(new_n8737));
  inv1 g08544(.a(new_n8737), .O(new_n8738));
  nor2 g08545(.a(new_n8690), .b(new_n8684), .O(new_n8739));
  inv1 g08546(.a(new_n8739), .O(new_n8740));
  nor2 g08547(.a(new_n8740), .b(new_n8738), .O(new_n8741));
  nor2 g08548(.a(new_n8739), .b(new_n8737), .O(new_n8742));
  nor2 g08549(.a(new_n8742), .b(new_n8741), .O(new_n8743));
  inv1 g08550(.a(new_n8743), .O(new_n8744));
  inv1 g08551(.a(new_n8472), .O(new_n8745));
  nor2 g08552(.a(new_n8745), .b(\a[54] ), .O(new_n8746));
  nor2 g08553(.a(new_n8476), .b(new_n2433), .O(new_n8747));
  inv1 g08554(.a(new_n8747), .O(new_n8748));
  nor2 g08555(.a(new_n8748), .b(new_n194), .O(new_n8749));
  nor2 g08556(.a(new_n8476), .b(new_n194), .O(new_n8750));
  nor2 g08557(.a(new_n8750), .b(\a[28] ), .O(new_n8751));
  nor2 g08558(.a(new_n8751), .b(new_n8749), .O(new_n8752));
  nor2 g08559(.a(new_n8752), .b(new_n8472), .O(new_n8753));
  nor2 g08560(.a(new_n8753), .b(new_n8746), .O(new_n8754));
  inv1 g08561(.a(new_n8754), .O(new_n8755));
  nor2 g08562(.a(new_n8599), .b(new_n8594), .O(new_n8756));
  inv1 g08563(.a(new_n8756), .O(new_n8757));
  nor2 g08564(.a(new_n8757), .b(new_n8755), .O(new_n8758));
  nor2 g08565(.a(new_n8756), .b(new_n8754), .O(new_n8759));
  nor2 g08566(.a(new_n8759), .b(new_n8758), .O(new_n8760));
  inv1 g08567(.a(new_n8760), .O(new_n8761));
  nor2 g08568(.a(new_n8761), .b(new_n8744), .O(new_n8762));
  nor2 g08569(.a(new_n8760), .b(new_n8743), .O(new_n8763));
  nor2 g08570(.a(new_n8763), .b(new_n8762), .O(new_n8764));
  inv1 g08571(.a(new_n8764), .O(new_n8765));
  nor2 g08572(.a(new_n8765), .b(new_n8736), .O(new_n8766));
  inv1 g08573(.a(new_n8736), .O(new_n8767));
  nor2 g08574(.a(new_n8764), .b(new_n8767), .O(new_n8768));
  nor2 g08575(.a(new_n8768), .b(new_n8766), .O(new_n8769));
  inv1 g08576(.a(new_n8769), .O(new_n8770));
  nor2 g08577(.a(new_n8666), .b(new_n8660), .O(new_n8771));
  nor2 g08578(.a(new_n8633), .b(new_n8627), .O(new_n8772));
  nor2 g08579(.a(new_n8772), .b(new_n8771), .O(new_n8773));
  inv1 g08580(.a(new_n8771), .O(new_n8774));
  inv1 g08581(.a(new_n8772), .O(new_n8775));
  nor2 g08582(.a(new_n8775), .b(new_n8774), .O(new_n8776));
  nor2 g08583(.a(new_n8776), .b(new_n8773), .O(new_n8777));
  nor2 g08584(.a(new_n8610), .b(new_n8604), .O(new_n8778));
  nor2 g08585(.a(new_n8778), .b(new_n8777), .O(new_n8779));
  inv1 g08586(.a(new_n8777), .O(new_n8780));
  inv1 g08587(.a(new_n8778), .O(new_n8781));
  nor2 g08588(.a(new_n8781), .b(new_n8780), .O(new_n8782));
  nor2 g08589(.a(new_n8782), .b(new_n8779), .O(new_n8783));
  inv1 g08590(.a(new_n8783), .O(new_n8784));
  nor2 g08591(.a(new_n8487), .b(new_n8463), .O(new_n8785));
  nor2 g08592(.a(new_n8785), .b(new_n8784), .O(new_n8786));
  inv1 g08593(.a(new_n8785), .O(new_n8787));
  nor2 g08594(.a(new_n8787), .b(new_n8783), .O(new_n8788));
  nor2 g08595(.a(new_n8788), .b(new_n8786), .O(new_n8789));
  inv1 g08596(.a(new_n8789), .O(new_n8790));
  nor2 g08597(.a(new_n8483), .b(new_n8479), .O(new_n8791));
  inv1 g08598(.a(new_n8791), .O(new_n8792));
  nor2 g08599(.a(new_n8648), .b(new_n8641), .O(new_n8793));
  nor2 g08600(.a(new_n8793), .b(new_n8792), .O(new_n8794));
  inv1 g08601(.a(new_n8793), .O(new_n8795));
  nor2 g08602(.a(new_n8795), .b(new_n8791), .O(new_n8796));
  nor2 g08603(.a(new_n8796), .b(new_n8794), .O(new_n8797));
  inv1 g08604(.a(new_n8797), .O(new_n8798));
  nor2 g08605(.a(new_n7294), .b(new_n229), .O(new_n8799));
  inv1 g08606(.a(new_n8799), .O(new_n8800));
  nor2 g08607(.a(new_n4093), .b(new_n1086), .O(new_n8801));
  nor2 g08608(.a(new_n3870), .b(new_n1199), .O(new_n8802));
  nor2 g08609(.a(new_n8802), .b(new_n8801), .O(new_n8803));
  nor2 g08610(.a(new_n4093), .b(new_n1199), .O(new_n8804));
  inv1 g08611(.a(new_n8804), .O(new_n8805));
  nor2 g08612(.a(new_n8805), .b(new_n8150), .O(new_n8806));
  nor2 g08613(.a(new_n8806), .b(new_n8803), .O(new_n8807));
  nor2 g08614(.a(new_n8807), .b(new_n8800), .O(new_n8808));
  inv1 g08615(.a(new_n8807), .O(new_n8809));
  nor2 g08616(.a(new_n8809), .b(new_n8799), .O(new_n8810));
  nor2 g08617(.a(new_n8810), .b(new_n8808), .O(new_n8811));
  nor2 g08618(.a(new_n8811), .b(new_n8798), .O(new_n8812));
  inv1 g08619(.a(new_n8811), .O(new_n8813));
  nor2 g08620(.a(new_n8813), .b(new_n8797), .O(new_n8814));
  nor2 g08621(.a(new_n8814), .b(new_n8812), .O(new_n8815));
  inv1 g08622(.a(new_n8815), .O(new_n8816));
  nor2 g08623(.a(new_n8816), .b(new_n8790), .O(new_n8817));
  nor2 g08624(.a(new_n8815), .b(new_n8789), .O(new_n8818));
  nor2 g08625(.a(new_n8818), .b(new_n8817), .O(new_n8819));
  inv1 g08626(.a(new_n8819), .O(new_n8820));
  nor2 g08627(.a(new_n8820), .b(new_n8770), .O(new_n8821));
  nor2 g08628(.a(new_n8819), .b(new_n8769), .O(new_n8822));
  nor2 g08629(.a(new_n8822), .b(new_n8821), .O(new_n8823));
  nor2 g08630(.a(new_n8823), .b(new_n8735), .O(new_n8824));
  inv1 g08631(.a(new_n8823), .O(new_n8825));
  nor2 g08632(.a(new_n8825), .b(new_n8734), .O(new_n8826));
  nor2 g08633(.a(new_n8826), .b(new_n8824), .O(new_n8827));
  nor2 g08634(.a(new_n8496), .b(new_n8491), .O(new_n8828));
  nor2 g08635(.a(new_n8461), .b(new_n8454), .O(new_n8829));
  nor2 g08636(.a(new_n8447), .b(new_n8441), .O(new_n8830));
  nor2 g08637(.a(new_n8830), .b(new_n8829), .O(new_n8831));
  inv1 g08638(.a(new_n8829), .O(new_n8832));
  inv1 g08639(.a(new_n8830), .O(new_n8833));
  nor2 g08640(.a(new_n8833), .b(new_n8832), .O(new_n8834));
  nor2 g08641(.a(new_n8834), .b(new_n8831), .O(new_n8835));
  nor2 g08642(.a(new_n8589), .b(new_n8584), .O(new_n8836));
  nor2 g08643(.a(new_n8836), .b(new_n8835), .O(new_n8837));
  inv1 g08644(.a(new_n8835), .O(new_n8838));
  inv1 g08645(.a(new_n8836), .O(new_n8839));
  nor2 g08646(.a(new_n8839), .b(new_n8838), .O(new_n8840));
  nor2 g08647(.a(new_n8840), .b(new_n8837), .O(new_n8841));
  inv1 g08648(.a(new_n8841), .O(new_n8842));
  nor2 g08649(.a(new_n8668), .b(new_n8650), .O(new_n8843));
  inv1 g08650(.a(new_n8843), .O(new_n8844));
  nor2 g08651(.a(new_n8619), .b(new_n8612), .O(new_n8845));
  inv1 g08652(.a(new_n8845), .O(new_n8846));
  nor2 g08653(.a(new_n8846), .b(new_n8844), .O(new_n8847));
  nor2 g08654(.a(new_n8845), .b(new_n8843), .O(new_n8848));
  nor2 g08655(.a(new_n8848), .b(new_n8847), .O(new_n8849));
  inv1 g08656(.a(new_n8849), .O(new_n8850));
  nor2 g08657(.a(new_n8850), .b(new_n8842), .O(new_n8851));
  nor2 g08658(.a(new_n8849), .b(new_n8841), .O(new_n8852));
  nor2 g08659(.a(new_n8852), .b(new_n8851), .O(new_n8853));
  inv1 g08660(.a(new_n8853), .O(new_n8854));
  nor2 g08661(.a(new_n8854), .b(new_n8828), .O(new_n8855));
  inv1 g08662(.a(new_n8828), .O(new_n8856));
  nor2 g08663(.a(new_n8853), .b(new_n8856), .O(new_n8857));
  nor2 g08664(.a(new_n8857), .b(new_n8855), .O(new_n8858));
  inv1 g08665(.a(new_n8858), .O(new_n8859));
  nor2 g08666(.a(new_n8523), .b(new_n8517), .O(new_n8860));
  inv1 g08667(.a(new_n8860), .O(new_n8861));
  nor2 g08668(.a(new_n4425), .b(new_n847), .O(new_n8862));
  inv1 g08669(.a(new_n8862), .O(new_n8863));
  nor2 g08670(.a(new_n6570), .b(new_n322), .O(new_n8864));
  nor2 g08671(.a(new_n6893), .b(new_n295), .O(new_n8865));
  nor2 g08672(.a(new_n8865), .b(new_n8864), .O(new_n8866));
  nor2 g08673(.a(new_n6893), .b(new_n322), .O(new_n8867));
  inv1 g08674(.a(new_n8867), .O(new_n8868));
  nor2 g08675(.a(new_n8868), .b(new_n8638), .O(new_n8869));
  nor2 g08676(.a(new_n8869), .b(new_n8866), .O(new_n8870));
  nor2 g08677(.a(new_n8870), .b(new_n8863), .O(new_n8871));
  inv1 g08678(.a(new_n8870), .O(new_n8872));
  nor2 g08679(.a(new_n8872), .b(new_n8862), .O(new_n8873));
  nor2 g08680(.a(new_n8873), .b(new_n8871), .O(new_n8874));
  inv1 g08681(.a(new_n8874), .O(new_n8875));
  nor2 g08682(.a(new_n5971), .b(new_n438), .O(new_n8876));
  nor2 g08683(.a(new_n5178), .b(new_n613), .O(new_n8877));
  nor2 g08684(.a(new_n5796), .b(new_n502), .O(new_n8878));
  nor2 g08685(.a(new_n8878), .b(new_n8877), .O(new_n8879));
  nor2 g08686(.a(new_n5796), .b(new_n613), .O(new_n8880));
  inv1 g08687(.a(new_n8880), .O(new_n8881));
  nor2 g08688(.a(new_n8881), .b(new_n8227), .O(new_n8882));
  nor2 g08689(.a(new_n8882), .b(new_n8879), .O(new_n8883));
  inv1 g08690(.a(new_n8883), .O(new_n8884));
  nor2 g08691(.a(new_n8884), .b(new_n8876), .O(new_n8885));
  inv1 g08692(.a(new_n8876), .O(new_n8886));
  nor2 g08693(.a(new_n8883), .b(new_n8886), .O(new_n8887));
  nor2 g08694(.a(new_n8887), .b(new_n8885), .O(new_n8888));
  nor2 g08695(.a(new_n2433), .b(new_n2184), .O(new_n8889));
  nor2 g08696(.a(new_n2506), .b(new_n2121), .O(new_n8890));
  nor2 g08697(.a(new_n8890), .b(new_n8889), .O(new_n8891));
  inv1 g08698(.a(new_n8889), .O(new_n8892));
  inv1 g08699(.a(new_n8890), .O(new_n8893));
  nor2 g08700(.a(new_n8893), .b(new_n8892), .O(new_n8894));
  nor2 g08701(.a(new_n8894), .b(new_n8891), .O(new_n8895));
  nor2 g08702(.a(new_n8895), .b(new_n8245), .O(new_n8896));
  inv1 g08703(.a(new_n8895), .O(new_n8897));
  nor2 g08704(.a(new_n8897), .b(new_n8244), .O(new_n8898));
  nor2 g08705(.a(new_n8898), .b(new_n8896), .O(new_n8899));
  nor2 g08706(.a(new_n8899), .b(new_n8888), .O(new_n8900));
  inv1 g08707(.a(new_n8888), .O(new_n8901));
  inv1 g08708(.a(new_n8899), .O(new_n8902));
  nor2 g08709(.a(new_n8902), .b(new_n8901), .O(new_n8903));
  nor2 g08710(.a(new_n8903), .b(new_n8900), .O(new_n8904));
  nor2 g08711(.a(new_n8904), .b(new_n8875), .O(new_n8905));
  inv1 g08712(.a(new_n8904), .O(new_n8906));
  nor2 g08713(.a(new_n8906), .b(new_n8874), .O(new_n8907));
  nor2 g08714(.a(new_n8907), .b(new_n8905), .O(new_n8908));
  nor2 g08715(.a(new_n8908), .b(new_n8861), .O(new_n8909));
  inv1 g08716(.a(new_n8908), .O(new_n8910));
  nor2 g08717(.a(new_n8910), .b(new_n8860), .O(new_n8911));
  nor2 g08718(.a(new_n8911), .b(new_n8909), .O(new_n8912));
  inv1 g08719(.a(new_n8912), .O(new_n8913));
  nor2 g08720(.a(new_n3057), .b(new_n1647), .O(new_n8914));
  inv1 g08721(.a(new_n8914), .O(new_n8915));
  nor2 g08722(.a(new_n2826), .b(new_n1736), .O(new_n8916));
  nor2 g08723(.a(new_n8916), .b(new_n8455), .O(new_n8917));
  nor2 g08724(.a(new_n2826), .b(new_n1903), .O(new_n8918));
  inv1 g08725(.a(new_n8918), .O(new_n8919));
  nor2 g08726(.a(new_n8919), .b(new_n8258), .O(new_n8920));
  nor2 g08727(.a(new_n8920), .b(new_n8917), .O(new_n8921));
  nor2 g08728(.a(new_n8921), .b(new_n8915), .O(new_n8922));
  inv1 g08729(.a(new_n8921), .O(new_n8923));
  nor2 g08730(.a(new_n8923), .b(new_n8914), .O(new_n8924));
  nor2 g08731(.a(new_n8924), .b(new_n8922), .O(new_n8925));
  inv1 g08732(.a(new_n8925), .O(new_n8926));
  nor2 g08733(.a(new_n3722), .b(new_n1297), .O(new_n8927));
  inv1 g08734(.a(new_n8927), .O(new_n8928));
  nor2 g08735(.a(new_n3533), .b(new_n1425), .O(new_n8929));
  nor2 g08736(.a(new_n8929), .b(new_n8442), .O(new_n8930));
  nor2 g08737(.a(new_n3533), .b(new_n1493), .O(new_n8931));
  inv1 g08738(.a(new_n8931), .O(new_n8932));
  nor2 g08739(.a(new_n8932), .b(new_n8125), .O(new_n8933));
  nor2 g08740(.a(new_n8933), .b(new_n8930), .O(new_n8934));
  nor2 g08741(.a(new_n8934), .b(new_n8928), .O(new_n8935));
  inv1 g08742(.a(new_n8934), .O(new_n8936));
  nor2 g08743(.a(new_n8936), .b(new_n8927), .O(new_n8937));
  nor2 g08744(.a(new_n8937), .b(new_n8935), .O(new_n8938));
  nor2 g08745(.a(new_n8170), .b(new_n196), .O(new_n8939));
  nor2 g08746(.a(new_n8939), .b(new_n8628), .O(new_n8940));
  inv1 g08747(.a(new_n8133), .O(new_n8941));
  nor2 g08748(.a(new_n8170), .b(new_n214), .O(new_n8942));
  inv1 g08749(.a(new_n8942), .O(new_n8943));
  nor2 g08750(.a(new_n8943), .b(new_n8941), .O(new_n8944));
  nor2 g08751(.a(new_n8944), .b(new_n8940), .O(new_n8945));
  inv1 g08752(.a(\a[55] ), .O(new_n8946));
  nor2 g08753(.a(new_n8946), .b(new_n198), .O(new_n8947));
  inv1 g08754(.a(new_n8947), .O(new_n8948));
  nor2 g08755(.a(new_n8948), .b(new_n8945), .O(new_n8949));
  inv1 g08756(.a(new_n8945), .O(new_n8950));
  nor2 g08757(.a(new_n8947), .b(new_n8950), .O(new_n8951));
  nor2 g08758(.a(new_n8951), .b(new_n8949), .O(new_n8952));
  nor2 g08759(.a(new_n8952), .b(new_n8938), .O(new_n8953));
  inv1 g08760(.a(new_n8938), .O(new_n8954));
  inv1 g08761(.a(new_n8952), .O(new_n8955));
  nor2 g08762(.a(new_n8955), .b(new_n8954), .O(new_n8956));
  nor2 g08763(.a(new_n8956), .b(new_n8953), .O(new_n8957));
  nor2 g08764(.a(new_n8957), .b(new_n8926), .O(new_n8958));
  inv1 g08765(.a(new_n8957), .O(new_n8959));
  nor2 g08766(.a(new_n8959), .b(new_n8925), .O(new_n8960));
  nor2 g08767(.a(new_n8960), .b(new_n8958), .O(new_n8961));
  inv1 g08768(.a(new_n8961), .O(new_n8962));
  nor2 g08769(.a(new_n8962), .b(new_n8913), .O(new_n8963));
  nor2 g08770(.a(new_n8961), .b(new_n8912), .O(new_n8964));
  nor2 g08771(.a(new_n8964), .b(new_n8963), .O(new_n8965));
  inv1 g08772(.a(new_n8965), .O(new_n8966));
  nor2 g08773(.a(new_n8966), .b(new_n8859), .O(new_n8967));
  nor2 g08774(.a(new_n8965), .b(new_n8858), .O(new_n8968));
  nor2 g08775(.a(new_n8968), .b(new_n8967), .O(new_n8969));
  nor2 g08776(.a(new_n8969), .b(new_n8827), .O(new_n8970));
  inv1 g08777(.a(new_n8827), .O(new_n8971));
  inv1 g08778(.a(new_n8969), .O(new_n8972));
  nor2 g08779(.a(new_n8972), .b(new_n8971), .O(new_n8973));
  nor2 g08780(.a(new_n8973), .b(new_n8970), .O(new_n8974));
  inv1 g08781(.a(new_n8974), .O(new_n8975));
  nor2 g08782(.a(new_n8714), .b(new_n8575), .O(new_n8976));
  nor2 g08783(.a(new_n8710), .b(new_n8705), .O(new_n8977));
  nor2 g08784(.a(new_n8570), .b(new_n8527), .O(new_n8978));
  nor2 g08785(.a(new_n8566), .b(new_n8563), .O(new_n8979));
  nor2 g08786(.a(new_n8557), .b(new_n8551), .O(new_n8980));
  inv1 g08787(.a(new_n8980), .O(new_n8981));
  nor2 g08788(.a(new_n8026), .b(new_n203), .O(new_n8982));
  nor2 g08789(.a(new_n6958), .b(new_n257), .O(new_n8983));
  nor2 g08790(.a(new_n4366), .b(new_n941), .O(new_n8984));
  nor2 g08791(.a(new_n8984), .b(new_n8983), .O(new_n8985));
  nor2 g08792(.a(new_n6958), .b(new_n941), .O(new_n8986));
  inv1 g08793(.a(new_n8986), .O(new_n8987));
  nor2 g08794(.a(new_n8987), .b(new_n5662), .O(new_n8988));
  nor2 g08795(.a(new_n8988), .b(new_n8985), .O(new_n8989));
  inv1 g08796(.a(new_n8989), .O(new_n8990));
  nor2 g08797(.a(new_n8990), .b(new_n8982), .O(new_n8991));
  inv1 g08798(.a(new_n8982), .O(new_n8992));
  nor2 g08799(.a(new_n8989), .b(new_n8992), .O(new_n8993));
  nor2 g08800(.a(new_n8993), .b(new_n8991), .O(new_n8994));
  nor2 g08801(.a(new_n4682), .b(new_n800), .O(new_n8995));
  inv1 g08802(.a(new_n8995), .O(new_n8996));
  nor2 g08803(.a(new_n6274), .b(new_n363), .O(new_n8997));
  nor2 g08804(.a(new_n8997), .b(new_n6510), .O(new_n8998));
  inv1 g08805(.a(new_n8997), .O(new_n8999));
  nor2 g08806(.a(new_n8999), .b(new_n6511), .O(new_n9000));
  nor2 g08807(.a(new_n9000), .b(new_n8998), .O(new_n9001));
  nor2 g08808(.a(new_n9001), .b(new_n8996), .O(new_n9002));
  inv1 g08809(.a(new_n9001), .O(new_n9003));
  nor2 g08810(.a(new_n9003), .b(new_n8995), .O(new_n9004));
  nor2 g08811(.a(new_n9004), .b(new_n9002), .O(new_n9005));
  nor2 g08812(.a(new_n9005), .b(new_n8994), .O(new_n9006));
  inv1 g08813(.a(new_n8994), .O(new_n9007));
  inv1 g08814(.a(new_n9005), .O(new_n9008));
  nor2 g08815(.a(new_n9008), .b(new_n9007), .O(new_n9009));
  nor2 g08816(.a(new_n9009), .b(new_n9006), .O(new_n9010));
  nor2 g08817(.a(new_n9010), .b(new_n8981), .O(new_n9011));
  inv1 g08818(.a(new_n9010), .O(new_n9012));
  nor2 g08819(.a(new_n9012), .b(new_n8980), .O(new_n9013));
  nor2 g08820(.a(new_n9013), .b(new_n9011), .O(new_n9014));
  inv1 g08821(.a(new_n9014), .O(new_n9015));
  nor2 g08822(.a(new_n8701), .b(new_n8698), .O(new_n9016));
  nor2 g08823(.a(new_n9016), .b(new_n9015), .O(new_n9017));
  inv1 g08824(.a(new_n9016), .O(new_n9018));
  nor2 g08825(.a(new_n9018), .b(new_n9014), .O(new_n9019));
  nor2 g08826(.a(new_n9019), .b(new_n9017), .O(new_n9020));
  inv1 g08827(.a(new_n9020), .O(new_n9021));
  nor2 g08828(.a(new_n9021), .b(new_n8979), .O(new_n9022));
  inv1 g08829(.a(new_n8979), .O(new_n9023));
  nor2 g08830(.a(new_n9020), .b(new_n9023), .O(new_n9024));
  nor2 g08831(.a(new_n9024), .b(new_n9022), .O(new_n9025));
  inv1 g08832(.a(new_n9025), .O(new_n9026));
  nor2 g08833(.a(new_n9026), .b(new_n8978), .O(new_n9027));
  inv1 g08834(.a(new_n8978), .O(new_n9028));
  nor2 g08835(.a(new_n9025), .b(new_n9028), .O(new_n9029));
  nor2 g08836(.a(new_n9029), .b(new_n9027), .O(new_n9030));
  inv1 g08837(.a(new_n9030), .O(new_n9031));
  nor2 g08838(.a(new_n9031), .b(new_n8977), .O(new_n9032));
  inv1 g08839(.a(new_n8977), .O(new_n9033));
  nor2 g08840(.a(new_n9030), .b(new_n9033), .O(new_n9034));
  nor2 g08841(.a(new_n9034), .b(new_n9032), .O(new_n9035));
  inv1 g08842(.a(new_n9035), .O(new_n9036));
  nor2 g08843(.a(new_n9036), .b(new_n8976), .O(new_n9037));
  inv1 g08844(.a(new_n8976), .O(new_n9038));
  nor2 g08845(.a(new_n9035), .b(new_n9038), .O(new_n9039));
  nor2 g08846(.a(new_n9039), .b(new_n9037), .O(new_n9040));
  inv1 g08847(.a(new_n9040), .O(new_n9041));
  nor2 g08848(.a(new_n9041), .b(new_n8975), .O(new_n9042));
  nor2 g08849(.a(new_n9040), .b(new_n8974), .O(new_n9043));
  nor2 g08850(.a(new_n9043), .b(new_n9042), .O(new_n9044));
  inv1 g08851(.a(new_n9044), .O(new_n9045));
  nor2 g08852(.a(new_n9045), .b(new_n8733), .O(new_n9046));
  inv1 g08853(.a(new_n8733), .O(new_n9047));
  nor2 g08854(.a(new_n9044), .b(new_n9047), .O(new_n9048));
  nor2 g08855(.a(new_n9048), .b(new_n9046), .O(new_n9049));
  inv1 g08856(.a(new_n9049), .O(new_n9050));
  nor2 g08857(.a(new_n8730), .b(new_n8724), .O(new_n9051));
  nor2 g08858(.a(new_n9051), .b(new_n9050), .O(new_n9052));
  inv1 g08859(.a(new_n9051), .O(new_n9053));
  nor2 g08860(.a(new_n9053), .b(new_n9049), .O(new_n9054));
  nor2 g08861(.a(new_n9054), .b(new_n9052), .O(new_n9055));
  inv1 g08862(.a(new_n9055), .O(\asquared[56] ));
  nor2 g08863(.a(new_n9042), .b(new_n9037), .O(new_n9057));
  nor2 g08864(.a(new_n4682), .b(new_n847), .O(new_n9058));
  inv1 g08865(.a(new_n9058), .O(new_n9059));
  nor2 g08866(.a(new_n8867), .b(new_n6142), .O(new_n9060));
  inv1 g08867(.a(new_n7048), .O(new_n9061));
  nor2 g08868(.a(new_n6893), .b(new_n800), .O(new_n9062));
  inv1 g08869(.a(new_n9062), .O(new_n9063));
  nor2 g08870(.a(new_n9063), .b(new_n9061), .O(new_n9064));
  nor2 g08871(.a(new_n9064), .b(new_n9060), .O(new_n9065));
  nor2 g08872(.a(new_n9065), .b(new_n9059), .O(new_n9066));
  inv1 g08873(.a(new_n9065), .O(new_n9067));
  nor2 g08874(.a(new_n9067), .b(new_n9058), .O(new_n9068));
  nor2 g08875(.a(new_n9068), .b(new_n9066), .O(new_n9069));
  inv1 g08876(.a(new_n9069), .O(new_n9070));
  nor2 g08877(.a(new_n5971), .b(new_n502), .O(new_n9071));
  inv1 g08878(.a(new_n9071), .O(new_n9072));
  nor2 g08879(.a(new_n5796), .b(new_n569), .O(new_n9073));
  nor2 g08880(.a(new_n9073), .b(new_n7627), .O(new_n9074));
  nor2 g08881(.a(new_n8881), .b(new_n8245), .O(new_n9075));
  nor2 g08882(.a(new_n9075), .b(new_n9074), .O(new_n9076));
  nor2 g08883(.a(new_n9076), .b(new_n9072), .O(new_n9077));
  inv1 g08884(.a(new_n9076), .O(new_n9078));
  nor2 g08885(.a(new_n9078), .b(new_n9071), .O(new_n9079));
  nor2 g08886(.a(new_n9079), .b(new_n9077), .O(new_n9080));
  nor2 g08887(.a(new_n7294), .b(new_n257), .O(new_n9081));
  inv1 g08888(.a(new_n9081), .O(new_n9082));
  nor2 g08889(.a(new_n6958), .b(new_n295), .O(new_n9083));
  nor2 g08890(.a(new_n4425), .b(new_n941), .O(new_n9084));
  nor2 g08891(.a(new_n9084), .b(new_n9083), .O(new_n9085));
  inv1 g08892(.a(new_n9083), .O(new_n9086));
  inv1 g08893(.a(new_n9084), .O(new_n9087));
  nor2 g08894(.a(new_n9087), .b(new_n9086), .O(new_n9088));
  nor2 g08895(.a(new_n9088), .b(new_n9085), .O(new_n9089));
  nor2 g08896(.a(new_n9089), .b(new_n9082), .O(new_n9090));
  inv1 g08897(.a(new_n9089), .O(new_n9091));
  nor2 g08898(.a(new_n9091), .b(new_n9081), .O(new_n9092));
  nor2 g08899(.a(new_n9092), .b(new_n9090), .O(new_n9093));
  nor2 g08900(.a(new_n9093), .b(new_n9080), .O(new_n9094));
  inv1 g08901(.a(new_n9080), .O(new_n9095));
  inv1 g08902(.a(new_n9093), .O(new_n9096));
  nor2 g08903(.a(new_n9096), .b(new_n9095), .O(new_n9097));
  nor2 g08904(.a(new_n9097), .b(new_n9094), .O(new_n9098));
  nor2 g08905(.a(new_n9098), .b(new_n9070), .O(new_n9099));
  inv1 g08906(.a(new_n9098), .O(new_n9100));
  nor2 g08907(.a(new_n9100), .b(new_n9069), .O(new_n9101));
  nor2 g08908(.a(new_n9101), .b(new_n9099), .O(new_n9102));
  inv1 g08909(.a(new_n9102), .O(new_n9103));
  nor2 g08910(.a(new_n6570), .b(new_n363), .O(new_n9104));
  inv1 g08911(.a(new_n9104), .O(new_n9105));
  nor2 g08912(.a(new_n5178), .b(new_n699), .O(new_n9106));
  nor2 g08913(.a(new_n6274), .b(new_n438), .O(new_n9107));
  nor2 g08914(.a(new_n9107), .b(new_n9106), .O(new_n9108));
  nor2 g08915(.a(new_n6274), .b(new_n699), .O(new_n9109));
  inv1 g08916(.a(new_n9109), .O(new_n9110));
  nor2 g08917(.a(new_n9110), .b(new_n7839), .O(new_n9111));
  nor2 g08918(.a(new_n9111), .b(new_n9108), .O(new_n9112));
  nor2 g08919(.a(new_n9112), .b(new_n9105), .O(new_n9113));
  inv1 g08920(.a(new_n9112), .O(new_n9114));
  nor2 g08921(.a(new_n9114), .b(new_n9104), .O(new_n9115));
  nor2 g08922(.a(new_n9115), .b(new_n9113), .O(new_n9116));
  inv1 g08923(.a(new_n9116), .O(new_n9117));
  nor2 g08924(.a(new_n3870), .b(new_n1297), .O(new_n9118));
  nor2 g08925(.a(new_n3231), .b(new_n1647), .O(new_n9119));
  nor2 g08926(.a(new_n9119), .b(new_n8931), .O(new_n9120));
  nor2 g08927(.a(new_n3533), .b(new_n1647), .O(new_n9121));
  inv1 g08928(.a(new_n9121), .O(new_n9122));
  nor2 g08929(.a(new_n9122), .b(new_n8443), .O(new_n9123));
  nor2 g08930(.a(new_n9123), .b(new_n9120), .O(new_n9124));
  inv1 g08931(.a(new_n9124), .O(new_n9125));
  nor2 g08932(.a(new_n9125), .b(new_n9118), .O(new_n9126));
  inv1 g08933(.a(new_n9118), .O(new_n9127));
  nor2 g08934(.a(new_n9124), .b(new_n9127), .O(new_n9128));
  nor2 g08935(.a(new_n9128), .b(new_n9126), .O(new_n9129));
  nor2 g08936(.a(new_n3057), .b(new_n1736), .O(new_n9130));
  inv1 g08937(.a(new_n9130), .O(new_n9131));
  nor2 g08938(.a(new_n2660), .b(new_n2121), .O(new_n9132));
  nor2 g08939(.a(new_n9132), .b(new_n8918), .O(new_n9133));
  nor2 g08940(.a(new_n2826), .b(new_n2121), .O(new_n9134));
  inv1 g08941(.a(new_n9134), .O(new_n9135));
  nor2 g08942(.a(new_n9135), .b(new_n8456), .O(new_n9136));
  nor2 g08943(.a(new_n9136), .b(new_n9133), .O(new_n9137));
  nor2 g08944(.a(new_n9137), .b(new_n9131), .O(new_n9138));
  inv1 g08945(.a(new_n9137), .O(new_n9139));
  nor2 g08946(.a(new_n9139), .b(new_n9130), .O(new_n9140));
  nor2 g08947(.a(new_n9140), .b(new_n9138), .O(new_n9141));
  nor2 g08948(.a(new_n9141), .b(new_n9129), .O(new_n9142));
  inv1 g08949(.a(new_n9129), .O(new_n9143));
  inv1 g08950(.a(new_n9141), .O(new_n9144));
  nor2 g08951(.a(new_n9144), .b(new_n9143), .O(new_n9145));
  nor2 g08952(.a(new_n9145), .b(new_n9142), .O(new_n9146));
  nor2 g08953(.a(new_n9146), .b(new_n9117), .O(new_n9147));
  inv1 g08954(.a(new_n9146), .O(new_n9148));
  nor2 g08955(.a(new_n9148), .b(new_n9116), .O(new_n9149));
  nor2 g08956(.a(new_n9149), .b(new_n9147), .O(new_n9150));
  inv1 g08957(.a(new_n9150), .O(new_n9151));
  nor2 g08958(.a(new_n9151), .b(new_n9103), .O(new_n9152));
  nor2 g08959(.a(new_n9150), .b(new_n9102), .O(new_n9153));
  nor2 g08960(.a(new_n9153), .b(new_n9152), .O(new_n9154));
  inv1 g08961(.a(new_n8749), .O(new_n9155));
  inv1 g08962(.a(\a[56] ), .O(new_n9156));
  nor2 g08963(.a(new_n9156), .b(new_n198), .O(new_n9157));
  nor2 g08964(.a(new_n8476), .b(new_n196), .O(new_n9158));
  nor2 g08965(.a(new_n9158), .b(new_n9157), .O(new_n9159));
  nor2 g08966(.a(new_n9156), .b(new_n196), .O(new_n9160));
  inv1 g08967(.a(new_n9160), .O(new_n9161));
  nor2 g08968(.a(new_n9161), .b(new_n8478), .O(new_n9162));
  nor2 g08969(.a(new_n9162), .b(new_n9159), .O(new_n9163));
  inv1 g08970(.a(new_n9163), .O(new_n9164));
  nor2 g08971(.a(new_n9164), .b(new_n9155), .O(new_n9165));
  nor2 g08972(.a(new_n9163), .b(new_n8749), .O(new_n9166));
  nor2 g08973(.a(new_n9166), .b(new_n9165), .O(new_n9167));
  inv1 g08974(.a(new_n9167), .O(new_n9168));
  nor2 g08975(.a(new_n8873), .b(new_n8866), .O(new_n9169));
  inv1 g08976(.a(new_n9169), .O(new_n9170));
  nor2 g08977(.a(new_n9170), .b(new_n9168), .O(new_n9171));
  nor2 g08978(.a(new_n9169), .b(new_n9167), .O(new_n9172));
  nor2 g08979(.a(new_n9172), .b(new_n9171), .O(new_n9173));
  inv1 g08980(.a(new_n9173), .O(new_n9174));
  nor2 g08981(.a(new_n8170), .b(new_n203), .O(new_n9175));
  inv1 g08982(.a(new_n9175), .O(new_n9176));
  nor2 g08983(.a(new_n8026), .b(new_n214), .O(new_n9177));
  nor2 g08984(.a(new_n9177), .b(new_n8804), .O(new_n9178));
  inv1 g08985(.a(new_n9177), .O(new_n9179));
  nor2 g08986(.a(new_n9179), .b(new_n8805), .O(new_n9180));
  nor2 g08987(.a(new_n9180), .b(new_n9178), .O(new_n9181));
  nor2 g08988(.a(new_n9181), .b(new_n9176), .O(new_n9182));
  inv1 g08989(.a(new_n9181), .O(new_n9183));
  nor2 g08990(.a(new_n9183), .b(new_n9175), .O(new_n9184));
  nor2 g08991(.a(new_n9184), .b(new_n9182), .O(new_n9185));
  nor2 g08992(.a(new_n9185), .b(new_n9174), .O(new_n9186));
  inv1 g08993(.a(new_n9185), .O(new_n9187));
  nor2 g08994(.a(new_n9187), .b(new_n9173), .O(new_n9188));
  nor2 g08995(.a(new_n9188), .b(new_n9186), .O(new_n9189));
  nor2 g08996(.a(new_n9189), .b(new_n9154), .O(new_n9190));
  inv1 g08997(.a(new_n9154), .O(new_n9191));
  inv1 g08998(.a(new_n9189), .O(new_n9192));
  nor2 g08999(.a(new_n9192), .b(new_n9191), .O(new_n9193));
  nor2 g09000(.a(new_n9193), .b(new_n9190), .O(new_n9194));
  inv1 g09001(.a(new_n9194), .O(new_n9195));
  nor2 g09002(.a(new_n9022), .b(new_n9017), .O(new_n9196));
  nor2 g09003(.a(new_n8937), .b(new_n8930), .O(new_n9197));
  nor2 g09004(.a(new_n8924), .b(new_n8917), .O(new_n9198));
  nor2 g09005(.a(new_n9198), .b(new_n9197), .O(new_n9199));
  inv1 g09006(.a(new_n9197), .O(new_n9200));
  inv1 g09007(.a(new_n9198), .O(new_n9201));
  nor2 g09008(.a(new_n9201), .b(new_n9200), .O(new_n9202));
  nor2 g09009(.a(new_n9202), .b(new_n9199), .O(new_n9203));
  nor2 g09010(.a(new_n8991), .b(new_n8985), .O(new_n9204));
  nor2 g09011(.a(new_n9204), .b(new_n9203), .O(new_n9205));
  inv1 g09012(.a(new_n9203), .O(new_n9206));
  inv1 g09013(.a(new_n9204), .O(new_n9207));
  nor2 g09014(.a(new_n9207), .b(new_n9206), .O(new_n9208));
  nor2 g09015(.a(new_n9208), .b(new_n9205), .O(new_n9209));
  inv1 g09016(.a(new_n9209), .O(new_n9210));
  nor2 g09017(.a(new_n2506), .b(new_n2184), .O(new_n9211));
  nor2 g09018(.a(new_n8946), .b(new_n194), .O(new_n9212));
  nor2 g09019(.a(new_n9212), .b(new_n9211), .O(new_n9213));
  inv1 g09020(.a(new_n9211), .O(new_n9214));
  inv1 g09021(.a(new_n9212), .O(new_n9215));
  nor2 g09022(.a(new_n9215), .b(new_n9214), .O(new_n9216));
  nor2 g09023(.a(new_n9216), .b(new_n9213), .O(new_n9217));
  inv1 g09024(.a(new_n9217), .O(new_n9218));
  nor2 g09025(.a(new_n8898), .b(new_n8891), .O(new_n9219));
  inv1 g09026(.a(new_n9219), .O(new_n9220));
  nor2 g09027(.a(new_n9220), .b(new_n9218), .O(new_n9221));
  nor2 g09028(.a(new_n9219), .b(new_n9217), .O(new_n9222));
  nor2 g09029(.a(new_n9222), .b(new_n9221), .O(new_n9223));
  inv1 g09030(.a(new_n9223), .O(new_n9224));
  nor2 g09031(.a(new_n8885), .b(new_n8879), .O(new_n9225));
  inv1 g09032(.a(new_n9225), .O(new_n9226));
  nor2 g09033(.a(new_n9226), .b(new_n9224), .O(new_n9227));
  nor2 g09034(.a(new_n9225), .b(new_n9223), .O(new_n9228));
  nor2 g09035(.a(new_n9228), .b(new_n9227), .O(new_n9229));
  inv1 g09036(.a(new_n9229), .O(new_n9230));
  nor2 g09037(.a(new_n8907), .b(new_n8900), .O(new_n9231));
  nor2 g09038(.a(new_n9231), .b(new_n9230), .O(new_n9232));
  inv1 g09039(.a(new_n9231), .O(new_n9233));
  nor2 g09040(.a(new_n9233), .b(new_n9229), .O(new_n9234));
  nor2 g09041(.a(new_n9234), .b(new_n9232), .O(new_n9235));
  inv1 g09042(.a(new_n9235), .O(new_n9236));
  nor2 g09043(.a(new_n9236), .b(new_n9210), .O(new_n9237));
  nor2 g09044(.a(new_n9235), .b(new_n9209), .O(new_n9238));
  nor2 g09045(.a(new_n9238), .b(new_n9237), .O(new_n9239));
  inv1 g09046(.a(new_n9239), .O(new_n9240));
  nor2 g09047(.a(new_n9240), .b(new_n9196), .O(new_n9241));
  inv1 g09048(.a(new_n9196), .O(new_n9242));
  nor2 g09049(.a(new_n9239), .b(new_n9242), .O(new_n9243));
  nor2 g09050(.a(new_n9243), .b(new_n9241), .O(new_n9244));
  inv1 g09051(.a(new_n9244), .O(new_n9245));
  nor2 g09052(.a(new_n9245), .b(new_n9195), .O(new_n9246));
  nor2 g09053(.a(new_n9244), .b(new_n9194), .O(new_n9247));
  nor2 g09054(.a(new_n9247), .b(new_n9246), .O(new_n9248));
  inv1 g09055(.a(new_n9248), .O(new_n9249));
  nor2 g09056(.a(new_n9032), .b(new_n9027), .O(new_n9250));
  nor2 g09057(.a(new_n8810), .b(new_n8803), .O(new_n9251));
  nor2 g09058(.a(new_n8951), .b(new_n8940), .O(new_n9252));
  nor2 g09059(.a(new_n9252), .b(new_n9251), .O(new_n9253));
  inv1 g09060(.a(new_n9251), .O(new_n9254));
  inv1 g09061(.a(new_n9252), .O(new_n9255));
  nor2 g09062(.a(new_n9255), .b(new_n9254), .O(new_n9256));
  nor2 g09063(.a(new_n9256), .b(new_n9253), .O(new_n9257));
  nor2 g09064(.a(new_n9004), .b(new_n8998), .O(new_n9258));
  nor2 g09065(.a(new_n9258), .b(new_n9257), .O(new_n9259));
  inv1 g09066(.a(new_n9257), .O(new_n9260));
  inv1 g09067(.a(new_n9258), .O(new_n9261));
  nor2 g09068(.a(new_n9261), .b(new_n9260), .O(new_n9262));
  nor2 g09069(.a(new_n9262), .b(new_n9259), .O(new_n9263));
  nor2 g09070(.a(new_n9013), .b(new_n9006), .O(new_n9264));
  inv1 g09071(.a(new_n9264), .O(new_n9265));
  nor2 g09072(.a(new_n9265), .b(new_n9263), .O(new_n9266));
  inv1 g09073(.a(new_n9263), .O(new_n9267));
  nor2 g09074(.a(new_n9264), .b(new_n9267), .O(new_n9268));
  nor2 g09075(.a(new_n9268), .b(new_n9266), .O(new_n9269));
  nor2 g09076(.a(new_n8762), .b(new_n8742), .O(new_n9270));
  inv1 g09077(.a(new_n9270), .O(new_n9271));
  nor2 g09078(.a(new_n9271), .b(new_n9269), .O(new_n9272));
  inv1 g09079(.a(new_n9269), .O(new_n9273));
  nor2 g09080(.a(new_n9270), .b(new_n9273), .O(new_n9274));
  nor2 g09081(.a(new_n9274), .b(new_n9272), .O(new_n9275));
  inv1 g09082(.a(new_n9275), .O(new_n9276));
  nor2 g09083(.a(new_n8840), .b(new_n8834), .O(new_n9277));
  inv1 g09084(.a(new_n9277), .O(new_n9278));
  nor2 g09085(.a(new_n8812), .b(new_n8796), .O(new_n9279));
  inv1 g09086(.a(new_n9279), .O(new_n9280));
  nor2 g09087(.a(new_n9280), .b(new_n9278), .O(new_n9281));
  nor2 g09088(.a(new_n9279), .b(new_n9277), .O(new_n9282));
  nor2 g09089(.a(new_n9282), .b(new_n9281), .O(new_n9283));
  nor2 g09090(.a(new_n8960), .b(new_n8953), .O(new_n9284));
  inv1 g09091(.a(new_n9284), .O(new_n9285));
  nor2 g09092(.a(new_n9285), .b(new_n9283), .O(new_n9286));
  inv1 g09093(.a(new_n9283), .O(new_n9287));
  nor2 g09094(.a(new_n9284), .b(new_n9287), .O(new_n9288));
  nor2 g09095(.a(new_n9288), .b(new_n9286), .O(new_n9289));
  inv1 g09096(.a(new_n9289), .O(new_n9290));
  nor2 g09097(.a(new_n8963), .b(new_n8911), .O(new_n9291));
  nor2 g09098(.a(new_n9291), .b(new_n9290), .O(new_n9292));
  inv1 g09099(.a(new_n9291), .O(new_n9293));
  nor2 g09100(.a(new_n9293), .b(new_n9289), .O(new_n9294));
  nor2 g09101(.a(new_n9294), .b(new_n9292), .O(new_n9295));
  inv1 g09102(.a(new_n9295), .O(new_n9296));
  nor2 g09103(.a(new_n9296), .b(new_n9276), .O(new_n9297));
  nor2 g09104(.a(new_n9295), .b(new_n9275), .O(new_n9298));
  nor2 g09105(.a(new_n9298), .b(new_n9297), .O(new_n9299));
  inv1 g09106(.a(new_n9299), .O(new_n9300));
  nor2 g09107(.a(new_n9300), .b(new_n9250), .O(new_n9301));
  inv1 g09108(.a(new_n9250), .O(new_n9302));
  nor2 g09109(.a(new_n9299), .b(new_n9302), .O(new_n9303));
  nor2 g09110(.a(new_n9303), .b(new_n9301), .O(new_n9304));
  inv1 g09111(.a(new_n9304), .O(new_n9305));
  nor2 g09112(.a(new_n9305), .b(new_n9249), .O(new_n9306));
  nor2 g09113(.a(new_n9304), .b(new_n9248), .O(new_n9307));
  nor2 g09114(.a(new_n9307), .b(new_n9306), .O(new_n9308));
  inv1 g09115(.a(new_n9308), .O(new_n9309));
  nor2 g09116(.a(new_n8782), .b(new_n8776), .O(new_n9310));
  inv1 g09117(.a(new_n9310), .O(new_n9311));
  nor2 g09118(.a(new_n8758), .b(new_n8746), .O(new_n9312));
  nor2 g09119(.a(new_n3722), .b(new_n1425), .O(new_n9313));
  inv1 g09120(.a(new_n9313), .O(new_n9314));
  nor2 g09121(.a(new_n7537), .b(new_n229), .O(new_n9315));
  nor2 g09122(.a(new_n4366), .b(new_n1086), .O(new_n9316));
  nor2 g09123(.a(new_n9316), .b(new_n9315), .O(new_n9317));
  nor2 g09124(.a(new_n7537), .b(new_n1086), .O(new_n9318));
  inv1 g09125(.a(new_n9318), .O(new_n9319));
  nor2 g09126(.a(new_n9319), .b(new_n5418), .O(new_n9320));
  nor2 g09127(.a(new_n9320), .b(new_n9317), .O(new_n9321));
  nor2 g09128(.a(new_n9321), .b(new_n9314), .O(new_n9322));
  inv1 g09129(.a(new_n9321), .O(new_n9323));
  nor2 g09130(.a(new_n9323), .b(new_n9313), .O(new_n9324));
  nor2 g09131(.a(new_n9324), .b(new_n9322), .O(new_n9325));
  nor2 g09132(.a(new_n9325), .b(new_n9312), .O(new_n9326));
  inv1 g09133(.a(new_n9312), .O(new_n9327));
  inv1 g09134(.a(new_n9325), .O(new_n9328));
  nor2 g09135(.a(new_n9328), .b(new_n9327), .O(new_n9329));
  nor2 g09136(.a(new_n9329), .b(new_n9326), .O(new_n9330));
  nor2 g09137(.a(new_n9330), .b(new_n9311), .O(new_n9331));
  inv1 g09138(.a(new_n9330), .O(new_n9332));
  nor2 g09139(.a(new_n9332), .b(new_n9310), .O(new_n9333));
  nor2 g09140(.a(new_n9333), .b(new_n9331), .O(new_n9334));
  inv1 g09141(.a(new_n9334), .O(new_n9335));
  nor2 g09142(.a(new_n8851), .b(new_n8848), .O(new_n9336));
  nor2 g09143(.a(new_n9336), .b(new_n9335), .O(new_n9337));
  inv1 g09144(.a(new_n9336), .O(new_n9338));
  nor2 g09145(.a(new_n9338), .b(new_n9334), .O(new_n9339));
  nor2 g09146(.a(new_n9339), .b(new_n9337), .O(new_n9340));
  nor2 g09147(.a(new_n8817), .b(new_n8786), .O(new_n9341));
  inv1 g09148(.a(new_n9341), .O(new_n9342));
  nor2 g09149(.a(new_n9342), .b(new_n9340), .O(new_n9343));
  inv1 g09150(.a(new_n9340), .O(new_n9344));
  nor2 g09151(.a(new_n9341), .b(new_n9344), .O(new_n9345));
  nor2 g09152(.a(new_n9345), .b(new_n9343), .O(new_n9346));
  nor2 g09153(.a(new_n8821), .b(new_n8766), .O(new_n9347));
  inv1 g09154(.a(new_n9347), .O(new_n9348));
  nor2 g09155(.a(new_n9348), .b(new_n9346), .O(new_n9349));
  inv1 g09156(.a(new_n9346), .O(new_n9350));
  nor2 g09157(.a(new_n9347), .b(new_n9350), .O(new_n9351));
  nor2 g09158(.a(new_n9351), .b(new_n9349), .O(new_n9352));
  nor2 g09159(.a(new_n8967), .b(new_n8855), .O(new_n9353));
  inv1 g09160(.a(new_n9353), .O(new_n9354));
  nor2 g09161(.a(new_n9354), .b(new_n9352), .O(new_n9355));
  inv1 g09162(.a(new_n9352), .O(new_n9356));
  nor2 g09163(.a(new_n9353), .b(new_n9356), .O(new_n9357));
  nor2 g09164(.a(new_n9357), .b(new_n9355), .O(new_n9358));
  inv1 g09165(.a(new_n9358), .O(new_n9359));
  nor2 g09166(.a(new_n8973), .b(new_n8826), .O(new_n9360));
  nor2 g09167(.a(new_n9360), .b(new_n9359), .O(new_n9361));
  inv1 g09168(.a(new_n9360), .O(new_n9362));
  nor2 g09169(.a(new_n9362), .b(new_n9358), .O(new_n9363));
  nor2 g09170(.a(new_n9363), .b(new_n9361), .O(new_n9364));
  inv1 g09171(.a(new_n9364), .O(new_n9365));
  nor2 g09172(.a(new_n9365), .b(new_n9309), .O(new_n9366));
  nor2 g09173(.a(new_n9364), .b(new_n9308), .O(new_n9367));
  nor2 g09174(.a(new_n9367), .b(new_n9366), .O(new_n9368));
  inv1 g09175(.a(new_n9368), .O(new_n9369));
  nor2 g09176(.a(new_n9369), .b(new_n9057), .O(new_n9370));
  inv1 g09177(.a(new_n9057), .O(new_n9371));
  nor2 g09178(.a(new_n9368), .b(new_n9371), .O(new_n9372));
  nor2 g09179(.a(new_n9372), .b(new_n9370), .O(new_n9373));
  inv1 g09180(.a(new_n9373), .O(new_n9374));
  nor2 g09181(.a(new_n9052), .b(new_n9048), .O(new_n9375));
  nor2 g09182(.a(new_n9375), .b(new_n9374), .O(new_n9376));
  inv1 g09183(.a(new_n9375), .O(new_n9377));
  nor2 g09184(.a(new_n9377), .b(new_n9373), .O(new_n9378));
  nor2 g09185(.a(new_n9378), .b(new_n9376), .O(new_n9379));
  inv1 g09186(.a(new_n9379), .O(\asquared[57] ));
  nor2 g09187(.a(new_n9366), .b(new_n9361), .O(new_n9381));
  nor2 g09188(.a(new_n9357), .b(new_n9351), .O(new_n9382));
  inv1 g09189(.a(new_n9382), .O(new_n9383));
  nor2 g09190(.a(new_n9227), .b(new_n9221), .O(new_n9384));
  inv1 g09191(.a(new_n9384), .O(new_n9385));
  nor2 g09192(.a(new_n9186), .b(new_n9171), .O(new_n9386));
  inv1 g09193(.a(new_n9386), .O(new_n9387));
  nor2 g09194(.a(new_n9387), .b(new_n9385), .O(new_n9388));
  nor2 g09195(.a(new_n9386), .b(new_n9384), .O(new_n9389));
  nor2 g09196(.a(new_n9389), .b(new_n9388), .O(new_n9390));
  nor2 g09197(.a(new_n9149), .b(new_n9142), .O(new_n9391));
  inv1 g09198(.a(new_n9391), .O(new_n9392));
  nor2 g09199(.a(new_n9392), .b(new_n9390), .O(new_n9393));
  inv1 g09200(.a(new_n9390), .O(new_n9394));
  nor2 g09201(.a(new_n9391), .b(new_n9394), .O(new_n9395));
  nor2 g09202(.a(new_n9395), .b(new_n9393), .O(new_n9396));
  inv1 g09203(.a(new_n9396), .O(new_n9397));
  nor2 g09204(.a(new_n9193), .b(new_n9152), .O(new_n9398));
  nor2 g09205(.a(new_n9398), .b(new_n9397), .O(new_n9399));
  inv1 g09206(.a(new_n9398), .O(new_n9400));
  nor2 g09207(.a(new_n9400), .b(new_n9396), .O(new_n9401));
  nor2 g09208(.a(new_n9401), .b(new_n9399), .O(new_n9402));
  inv1 g09209(.a(new_n9402), .O(new_n9403));
  nor2 g09210(.a(new_n9068), .b(new_n9060), .O(new_n9404));
  nor2 g09211(.a(new_n9140), .b(new_n9133), .O(new_n9405));
  nor2 g09212(.a(new_n9405), .b(new_n9404), .O(new_n9406));
  inv1 g09213(.a(new_n9404), .O(new_n9407));
  inv1 g09214(.a(new_n9405), .O(new_n9408));
  nor2 g09215(.a(new_n9408), .b(new_n9407), .O(new_n9409));
  nor2 g09216(.a(new_n9409), .b(new_n9406), .O(new_n9410));
  nor2 g09217(.a(new_n9092), .b(new_n9085), .O(new_n9411));
  nor2 g09218(.a(new_n9411), .b(new_n9410), .O(new_n9412));
  inv1 g09219(.a(new_n9410), .O(new_n9413));
  inv1 g09220(.a(new_n9411), .O(new_n9414));
  nor2 g09221(.a(new_n9414), .b(new_n9413), .O(new_n9415));
  nor2 g09222(.a(new_n9415), .b(new_n9412), .O(new_n9416));
  inv1 g09223(.a(new_n9416), .O(new_n9417));
  nor2 g09224(.a(new_n9184), .b(new_n9178), .O(new_n9418));
  nor2 g09225(.a(new_n9126), .b(new_n9120), .O(new_n9419));
  nor2 g09226(.a(new_n9419), .b(new_n9418), .O(new_n9420));
  inv1 g09227(.a(new_n9418), .O(new_n9421));
  inv1 g09228(.a(new_n9419), .O(new_n9422));
  nor2 g09229(.a(new_n9422), .b(new_n9421), .O(new_n9423));
  nor2 g09230(.a(new_n9423), .b(new_n9420), .O(new_n9424));
  nor2 g09231(.a(new_n9165), .b(new_n9162), .O(new_n9425));
  inv1 g09232(.a(new_n9425), .O(new_n9426));
  nor2 g09233(.a(new_n9426), .b(new_n9424), .O(new_n9427));
  inv1 g09234(.a(new_n9424), .O(new_n9428));
  nor2 g09235(.a(new_n9425), .b(new_n9428), .O(new_n9429));
  nor2 g09236(.a(new_n9429), .b(new_n9427), .O(new_n9430));
  inv1 g09237(.a(new_n9430), .O(new_n9431));
  nor2 g09238(.a(new_n9431), .b(new_n9417), .O(new_n9432));
  nor2 g09239(.a(new_n9430), .b(new_n9416), .O(new_n9433));
  nor2 g09240(.a(new_n9433), .b(new_n9432), .O(new_n9434));
  inv1 g09241(.a(new_n9434), .O(new_n9435));
  nor2 g09242(.a(new_n9101), .b(new_n9094), .O(new_n9436));
  nor2 g09243(.a(new_n9436), .b(new_n9435), .O(new_n9437));
  inv1 g09244(.a(new_n9436), .O(new_n9438));
  nor2 g09245(.a(new_n9438), .b(new_n9434), .O(new_n9439));
  nor2 g09246(.a(new_n9439), .b(new_n9437), .O(new_n9440));
  inv1 g09247(.a(new_n9440), .O(new_n9441));
  nor2 g09248(.a(new_n9441), .b(new_n9403), .O(new_n9442));
  nor2 g09249(.a(new_n9440), .b(new_n9402), .O(new_n9443));
  nor2 g09250(.a(new_n9443), .b(new_n9442), .O(new_n9444));
  nor2 g09251(.a(new_n9444), .b(new_n9383), .O(new_n9445));
  inv1 g09252(.a(new_n9444), .O(new_n9446));
  nor2 g09253(.a(new_n9446), .b(new_n9382), .O(new_n9447));
  nor2 g09254(.a(new_n9447), .b(new_n9445), .O(new_n9448));
  inv1 g09255(.a(new_n9448), .O(new_n9449));
  nor2 g09256(.a(new_n9288), .b(new_n9282), .O(new_n9450));
  nor2 g09257(.a(new_n5178), .b(new_n800), .O(new_n9451));
  inv1 g09258(.a(new_n9451), .O(new_n9452));
  nor2 g09259(.a(new_n6893), .b(new_n363), .O(new_n9453));
  nor2 g09260(.a(new_n6570), .b(new_n438), .O(new_n9454));
  nor2 g09261(.a(new_n9454), .b(new_n9453), .O(new_n9455));
  nor2 g09262(.a(new_n6893), .b(new_n438), .O(new_n9456));
  inv1 g09263(.a(new_n9456), .O(new_n9457));
  nor2 g09264(.a(new_n9457), .b(new_n9105), .O(new_n9458));
  nor2 g09265(.a(new_n9458), .b(new_n9455), .O(new_n9459));
  nor2 g09266(.a(new_n9459), .b(new_n9452), .O(new_n9460));
  inv1 g09267(.a(new_n9459), .O(new_n9461));
  nor2 g09268(.a(new_n9461), .b(new_n9451), .O(new_n9462));
  nor2 g09269(.a(new_n9462), .b(new_n9460), .O(new_n9463));
  inv1 g09270(.a(new_n9463), .O(new_n9464));
  nor2 g09271(.a(new_n8476), .b(new_n203), .O(new_n9465));
  nor2 g09272(.a(new_n8946), .b(new_n196), .O(new_n9466));
  nor2 g09273(.a(new_n9466), .b(new_n8942), .O(new_n9467));
  inv1 g09274(.a(new_n8939), .O(new_n9468));
  nor2 g09275(.a(new_n8946), .b(new_n214), .O(new_n9469));
  inv1 g09276(.a(new_n9469), .O(new_n9470));
  nor2 g09277(.a(new_n9470), .b(new_n9468), .O(new_n9471));
  nor2 g09278(.a(new_n9471), .b(new_n9467), .O(new_n9472));
  inv1 g09279(.a(new_n9472), .O(new_n9473));
  nor2 g09280(.a(new_n9473), .b(new_n9465), .O(new_n9474));
  inv1 g09281(.a(new_n9465), .O(new_n9475));
  nor2 g09282(.a(new_n9472), .b(new_n9475), .O(new_n9476));
  nor2 g09283(.a(new_n9476), .b(new_n9474), .O(new_n9477));
  nor2 g09284(.a(new_n8026), .b(new_n229), .O(new_n9478));
  inv1 g09285(.a(new_n9478), .O(new_n9479));
  nor2 g09286(.a(new_n4366), .b(new_n1199), .O(new_n9480));
  nor2 g09287(.a(new_n4093), .b(new_n1297), .O(new_n9481));
  nor2 g09288(.a(new_n9481), .b(new_n9480), .O(new_n9482));
  nor2 g09289(.a(new_n4366), .b(new_n1297), .O(new_n9483));
  inv1 g09290(.a(new_n9483), .O(new_n9484));
  nor2 g09291(.a(new_n9484), .b(new_n8805), .O(new_n9485));
  nor2 g09292(.a(new_n9485), .b(new_n9482), .O(new_n9486));
  nor2 g09293(.a(new_n9486), .b(new_n9479), .O(new_n9487));
  inv1 g09294(.a(new_n9486), .O(new_n9488));
  nor2 g09295(.a(new_n9488), .b(new_n9478), .O(new_n9489));
  nor2 g09296(.a(new_n9489), .b(new_n9487), .O(new_n9490));
  nor2 g09297(.a(new_n9490), .b(new_n9477), .O(new_n9491));
  inv1 g09298(.a(new_n9477), .O(new_n9492));
  inv1 g09299(.a(new_n9490), .O(new_n9493));
  nor2 g09300(.a(new_n9493), .b(new_n9492), .O(new_n9494));
  nor2 g09301(.a(new_n9494), .b(new_n9491), .O(new_n9495));
  nor2 g09302(.a(new_n9495), .b(new_n9464), .O(new_n9496));
  inv1 g09303(.a(new_n9495), .O(new_n9497));
  nor2 g09304(.a(new_n9497), .b(new_n9463), .O(new_n9498));
  nor2 g09305(.a(new_n9498), .b(new_n9496), .O(new_n9499));
  nor2 g09306(.a(new_n4425), .b(new_n1086), .O(new_n9500));
  inv1 g09307(.a(new_n9500), .O(new_n9501));
  nor2 g09308(.a(new_n7537), .b(new_n257), .O(new_n9502));
  nor2 g09309(.a(new_n4682), .b(new_n941), .O(new_n9503));
  nor2 g09310(.a(new_n9503), .b(new_n9502), .O(new_n9504));
  nor2 g09311(.a(new_n7537), .b(new_n941), .O(new_n9505));
  inv1 g09312(.a(new_n9505), .O(new_n9506));
  nor2 g09313(.a(new_n9506), .b(new_n6155), .O(new_n9507));
  nor2 g09314(.a(new_n9507), .b(new_n9504), .O(new_n9508));
  nor2 g09315(.a(new_n9508), .b(new_n9501), .O(new_n9509));
  inv1 g09316(.a(new_n9508), .O(new_n9510));
  nor2 g09317(.a(new_n9510), .b(new_n9500), .O(new_n9511));
  nor2 g09318(.a(new_n9511), .b(new_n9509), .O(new_n9512));
  inv1 g09319(.a(new_n9512), .O(new_n9513));
  nor2 g09320(.a(new_n6274), .b(new_n502), .O(new_n9514));
  nor2 g09321(.a(new_n9514), .b(new_n8880), .O(new_n9515));
  inv1 g09322(.a(new_n8878), .O(new_n9516));
  nor2 g09323(.a(new_n6274), .b(new_n613), .O(new_n9517));
  inv1 g09324(.a(new_n9517), .O(new_n9518));
  nor2 g09325(.a(new_n9518), .b(new_n9516), .O(new_n9519));
  nor2 g09326(.a(new_n9519), .b(new_n9515), .O(new_n9520));
  inv1 g09327(.a(new_n9520), .O(new_n9521));
  nor2 g09328(.a(new_n9521), .b(new_n7038), .O(new_n9522));
  nor2 g09329(.a(new_n9520), .b(new_n7039), .O(new_n9523));
  nor2 g09330(.a(new_n9523), .b(new_n9522), .O(new_n9524));
  nor2 g09331(.a(new_n5971), .b(new_n569), .O(new_n9525));
  inv1 g09332(.a(new_n9525), .O(new_n9526));
  nor2 g09333(.a(new_n2506), .b(new_n2433), .O(new_n9527));
  nor2 g09334(.a(new_n2660), .b(new_n2184), .O(new_n9528));
  nor2 g09335(.a(new_n9528), .b(new_n9527), .O(new_n9529));
  nor2 g09336(.a(new_n2660), .b(new_n2433), .O(new_n9530));
  inv1 g09337(.a(new_n9530), .O(new_n9531));
  nor2 g09338(.a(new_n9531), .b(new_n9214), .O(new_n9532));
  nor2 g09339(.a(new_n9532), .b(new_n9529), .O(new_n9533));
  nor2 g09340(.a(new_n9533), .b(new_n9526), .O(new_n9534));
  inv1 g09341(.a(new_n9533), .O(new_n9535));
  nor2 g09342(.a(new_n9535), .b(new_n9525), .O(new_n9536));
  nor2 g09343(.a(new_n9536), .b(new_n9534), .O(new_n9537));
  nor2 g09344(.a(new_n9537), .b(new_n9524), .O(new_n9538));
  inv1 g09345(.a(new_n9524), .O(new_n9539));
  inv1 g09346(.a(new_n9537), .O(new_n9540));
  nor2 g09347(.a(new_n9540), .b(new_n9539), .O(new_n9541));
  nor2 g09348(.a(new_n9541), .b(new_n9538), .O(new_n9542));
  nor2 g09349(.a(new_n9542), .b(new_n9513), .O(new_n9543));
  inv1 g09350(.a(new_n9542), .O(new_n9544));
  nor2 g09351(.a(new_n9544), .b(new_n9512), .O(new_n9545));
  nor2 g09352(.a(new_n9545), .b(new_n9543), .O(new_n9546));
  nor2 g09353(.a(new_n9546), .b(new_n9499), .O(new_n9547));
  inv1 g09354(.a(new_n9499), .O(new_n9548));
  inv1 g09355(.a(new_n9546), .O(new_n9549));
  nor2 g09356(.a(new_n9549), .b(new_n9548), .O(new_n9550));
  nor2 g09357(.a(new_n9550), .b(new_n9547), .O(new_n9551));
  inv1 g09358(.a(new_n9551), .O(new_n9552));
  nor2 g09359(.a(new_n9552), .b(new_n9450), .O(new_n9553));
  inv1 g09360(.a(new_n9450), .O(new_n9554));
  nor2 g09361(.a(new_n9551), .b(new_n9554), .O(new_n9555));
  nor2 g09362(.a(new_n9555), .b(new_n9553), .O(new_n9556));
  inv1 g09363(.a(new_n9556), .O(new_n9557));
  nor2 g09364(.a(new_n9345), .b(new_n9337), .O(new_n9558));
  nor2 g09365(.a(new_n9324), .b(new_n9317), .O(new_n9559));
  nor2 g09366(.a(new_n9115), .b(new_n9108), .O(new_n9560));
  nor2 g09367(.a(new_n9560), .b(new_n9559), .O(new_n9561));
  inv1 g09368(.a(new_n9559), .O(new_n9562));
  inv1 g09369(.a(new_n9560), .O(new_n9563));
  nor2 g09370(.a(new_n9563), .b(new_n9562), .O(new_n9564));
  nor2 g09371(.a(new_n9564), .b(new_n9561), .O(new_n9565));
  nor2 g09372(.a(new_n9079), .b(new_n9074), .O(new_n9566));
  nor2 g09373(.a(new_n9566), .b(new_n9565), .O(new_n9567));
  inv1 g09374(.a(new_n9565), .O(new_n9568));
  inv1 g09375(.a(new_n9566), .O(new_n9569));
  nor2 g09376(.a(new_n9569), .b(new_n9568), .O(new_n9570));
  nor2 g09377(.a(new_n9570), .b(new_n9567), .O(new_n9571));
  nor2 g09378(.a(new_n9333), .b(new_n9326), .O(new_n9572));
  inv1 g09379(.a(new_n9572), .O(new_n9573));
  nor2 g09380(.a(new_n9573), .b(new_n9571), .O(new_n9574));
  inv1 g09381(.a(new_n9571), .O(new_n9575));
  nor2 g09382(.a(new_n9572), .b(new_n9575), .O(new_n9576));
  nor2 g09383(.a(new_n9576), .b(new_n9574), .O(new_n9577));
  inv1 g09384(.a(new_n9577), .O(new_n9578));
  nor2 g09385(.a(new_n3231), .b(new_n1736), .O(new_n9579));
  inv1 g09386(.a(new_n9579), .O(new_n9580));
  nor2 g09387(.a(new_n3057), .b(new_n1903), .O(new_n9581));
  nor2 g09388(.a(new_n9581), .b(new_n9134), .O(new_n9582));
  nor2 g09389(.a(new_n3057), .b(new_n2121), .O(new_n9583));
  inv1 g09390(.a(new_n9583), .O(new_n9584));
  nor2 g09391(.a(new_n9584), .b(new_n8919), .O(new_n9585));
  nor2 g09392(.a(new_n9585), .b(new_n9582), .O(new_n9586));
  nor2 g09393(.a(new_n9586), .b(new_n9580), .O(new_n9587));
  inv1 g09394(.a(new_n9586), .O(new_n9588));
  nor2 g09395(.a(new_n9588), .b(new_n9579), .O(new_n9589));
  nor2 g09396(.a(new_n9589), .b(new_n9587), .O(new_n9590));
  inv1 g09397(.a(new_n9590), .O(new_n9591));
  nor2 g09398(.a(new_n7294), .b(new_n295), .O(new_n9592));
  nor2 g09399(.a(new_n6958), .b(new_n322), .O(new_n9593));
  nor2 g09400(.a(new_n4954), .b(new_n847), .O(new_n9594));
  nor2 g09401(.a(new_n9594), .b(new_n9593), .O(new_n9595));
  nor2 g09402(.a(new_n6958), .b(new_n847), .O(new_n9596));
  inv1 g09403(.a(new_n9596), .O(new_n9597));
  nor2 g09404(.a(new_n9597), .b(new_n9061), .O(new_n9598));
  nor2 g09405(.a(new_n9598), .b(new_n9595), .O(new_n9599));
  inv1 g09406(.a(new_n9599), .O(new_n9600));
  nor2 g09407(.a(new_n9600), .b(new_n9592), .O(new_n9601));
  inv1 g09408(.a(new_n9592), .O(new_n9602));
  nor2 g09409(.a(new_n9599), .b(new_n9602), .O(new_n9603));
  nor2 g09410(.a(new_n9603), .b(new_n9601), .O(new_n9604));
  nor2 g09411(.a(new_n3870), .b(new_n1425), .O(new_n9605));
  inv1 g09412(.a(new_n9605), .O(new_n9606));
  nor2 g09413(.a(new_n3722), .b(new_n1493), .O(new_n9607));
  nor2 g09414(.a(new_n9607), .b(new_n9121), .O(new_n9608));
  nor2 g09415(.a(new_n3722), .b(new_n1647), .O(new_n9609));
  inv1 g09416(.a(new_n9609), .O(new_n9610));
  nor2 g09417(.a(new_n9610), .b(new_n8932), .O(new_n9611));
  nor2 g09418(.a(new_n9611), .b(new_n9608), .O(new_n9612));
  nor2 g09419(.a(new_n9612), .b(new_n9606), .O(new_n9613));
  inv1 g09420(.a(new_n9612), .O(new_n9614));
  nor2 g09421(.a(new_n9614), .b(new_n9605), .O(new_n9615));
  nor2 g09422(.a(new_n9615), .b(new_n9613), .O(new_n9616));
  nor2 g09423(.a(new_n9616), .b(new_n9604), .O(new_n9617));
  inv1 g09424(.a(new_n9604), .O(new_n9618));
  inv1 g09425(.a(new_n9616), .O(new_n9619));
  nor2 g09426(.a(new_n9619), .b(new_n9618), .O(new_n9620));
  nor2 g09427(.a(new_n9620), .b(new_n9617), .O(new_n9621));
  nor2 g09428(.a(new_n9621), .b(new_n9591), .O(new_n9622));
  inv1 g09429(.a(new_n9621), .O(new_n9623));
  nor2 g09430(.a(new_n9623), .b(new_n9590), .O(new_n9624));
  nor2 g09431(.a(new_n9624), .b(new_n9622), .O(new_n9625));
  inv1 g09432(.a(new_n9625), .O(new_n9626));
  nor2 g09433(.a(new_n9626), .b(new_n9578), .O(new_n9627));
  nor2 g09434(.a(new_n9625), .b(new_n9577), .O(new_n9628));
  nor2 g09435(.a(new_n9628), .b(new_n9627), .O(new_n9629));
  inv1 g09436(.a(new_n9629), .O(new_n9630));
  nor2 g09437(.a(new_n9630), .b(new_n9558), .O(new_n9631));
  inv1 g09438(.a(new_n9558), .O(new_n9632));
  nor2 g09439(.a(new_n9629), .b(new_n9632), .O(new_n9633));
  nor2 g09440(.a(new_n9633), .b(new_n9631), .O(new_n9634));
  inv1 g09441(.a(new_n9634), .O(new_n9635));
  nor2 g09442(.a(new_n9635), .b(new_n9557), .O(new_n9636));
  nor2 g09443(.a(new_n9634), .b(new_n9556), .O(new_n9637));
  nor2 g09444(.a(new_n9637), .b(new_n9636), .O(new_n9638));
  inv1 g09445(.a(new_n9638), .O(new_n9639));
  nor2 g09446(.a(new_n9639), .b(new_n9449), .O(new_n9640));
  nor2 g09447(.a(new_n9638), .b(new_n9448), .O(new_n9641));
  nor2 g09448(.a(new_n9641), .b(new_n9640), .O(new_n9642));
  inv1 g09449(.a(new_n9642), .O(new_n9643));
  nor2 g09450(.a(new_n9306), .b(new_n9301), .O(new_n9644));
  nor2 g09451(.a(new_n9246), .b(new_n9241), .O(new_n9645));
  nor2 g09452(.a(new_n9297), .b(new_n9292), .O(new_n9646));
  nor2 g09453(.a(new_n9274), .b(new_n9268), .O(new_n9647));
  inv1 g09454(.a(new_n9647), .O(new_n9648));
  nor2 g09455(.a(new_n9237), .b(new_n9232), .O(new_n9649));
  inv1 g09456(.a(new_n9649), .O(new_n9650));
  nor2 g09457(.a(new_n9650), .b(new_n9648), .O(new_n9651));
  nor2 g09458(.a(new_n9649), .b(new_n9647), .O(new_n9652));
  nor2 g09459(.a(new_n9652), .b(new_n9651), .O(new_n9653));
  inv1 g09460(.a(new_n9653), .O(new_n9654));
  nor2 g09461(.a(new_n9208), .b(new_n9202), .O(new_n9655));
  inv1 g09462(.a(new_n9655), .O(new_n9656));
  inv1 g09463(.a(new_n9216), .O(new_n9657));
  inv1 g09464(.a(\a[57] ), .O(new_n9658));
  nor2 g09465(.a(new_n9658), .b(new_n198), .O(new_n9659));
  inv1 g09466(.a(new_n9659), .O(new_n9660));
  nor2 g09467(.a(new_n9660), .b(new_n9657), .O(new_n9661));
  nor2 g09468(.a(new_n9659), .b(new_n9216), .O(new_n9662));
  nor2 g09469(.a(new_n9662), .b(new_n9661), .O(new_n9663));
  inv1 g09470(.a(new_n9663), .O(new_n9664));
  nor2 g09471(.a(new_n9156), .b(new_n194), .O(new_n9665));
  inv1 g09472(.a(new_n9665), .O(new_n9666));
  nor2 g09473(.a(new_n9666), .b(new_n2506), .O(new_n9667));
  nor2 g09474(.a(new_n9665), .b(\a[29] ), .O(new_n9668));
  nor2 g09475(.a(new_n9668), .b(new_n9667), .O(new_n9669));
  inv1 g09476(.a(new_n9669), .O(new_n9670));
  nor2 g09477(.a(new_n9670), .b(new_n9664), .O(new_n9671));
  nor2 g09478(.a(new_n9669), .b(new_n9663), .O(new_n9672));
  nor2 g09479(.a(new_n9672), .b(new_n9671), .O(new_n9673));
  nor2 g09480(.a(new_n9673), .b(new_n9656), .O(new_n9674));
  inv1 g09481(.a(new_n9673), .O(new_n9675));
  nor2 g09482(.a(new_n9675), .b(new_n9655), .O(new_n9676));
  nor2 g09483(.a(new_n9676), .b(new_n9674), .O(new_n9677));
  nor2 g09484(.a(new_n9262), .b(new_n9256), .O(new_n9678));
  inv1 g09485(.a(new_n9678), .O(new_n9679));
  nor2 g09486(.a(new_n9679), .b(new_n9677), .O(new_n9680));
  inv1 g09487(.a(new_n9677), .O(new_n9681));
  nor2 g09488(.a(new_n9678), .b(new_n9681), .O(new_n9682));
  nor2 g09489(.a(new_n9682), .b(new_n9680), .O(new_n9683));
  inv1 g09490(.a(new_n9683), .O(new_n9684));
  nor2 g09491(.a(new_n9684), .b(new_n9654), .O(new_n9685));
  nor2 g09492(.a(new_n9683), .b(new_n9653), .O(new_n9686));
  nor2 g09493(.a(new_n9686), .b(new_n9685), .O(new_n9687));
  inv1 g09494(.a(new_n9687), .O(new_n9688));
  nor2 g09495(.a(new_n9688), .b(new_n9646), .O(new_n9689));
  inv1 g09496(.a(new_n9646), .O(new_n9690));
  nor2 g09497(.a(new_n9687), .b(new_n9690), .O(new_n9691));
  nor2 g09498(.a(new_n9691), .b(new_n9689), .O(new_n9692));
  inv1 g09499(.a(new_n9692), .O(new_n9693));
  nor2 g09500(.a(new_n9693), .b(new_n9645), .O(new_n9694));
  inv1 g09501(.a(new_n9645), .O(new_n9695));
  nor2 g09502(.a(new_n9692), .b(new_n9695), .O(new_n9696));
  nor2 g09503(.a(new_n9696), .b(new_n9694), .O(new_n9697));
  inv1 g09504(.a(new_n9697), .O(new_n9698));
  nor2 g09505(.a(new_n9698), .b(new_n9644), .O(new_n9699));
  inv1 g09506(.a(new_n9644), .O(new_n9700));
  nor2 g09507(.a(new_n9697), .b(new_n9700), .O(new_n9701));
  nor2 g09508(.a(new_n9701), .b(new_n9699), .O(new_n9702));
  inv1 g09509(.a(new_n9702), .O(new_n9703));
  nor2 g09510(.a(new_n9703), .b(new_n9643), .O(new_n9704));
  nor2 g09511(.a(new_n9702), .b(new_n9642), .O(new_n9705));
  nor2 g09512(.a(new_n9705), .b(new_n9704), .O(new_n9706));
  inv1 g09513(.a(new_n9706), .O(new_n9707));
  nor2 g09514(.a(new_n9707), .b(new_n9381), .O(new_n9708));
  inv1 g09515(.a(new_n9381), .O(new_n9709));
  nor2 g09516(.a(new_n9706), .b(new_n9709), .O(new_n9710));
  nor2 g09517(.a(new_n9710), .b(new_n9708), .O(new_n9711));
  inv1 g09518(.a(new_n9711), .O(new_n9712));
  nor2 g09519(.a(new_n9376), .b(new_n9372), .O(new_n9713));
  nor2 g09520(.a(new_n9713), .b(new_n9712), .O(new_n9714));
  inv1 g09521(.a(new_n9713), .O(new_n9715));
  nor2 g09522(.a(new_n9715), .b(new_n9711), .O(new_n9716));
  nor2 g09523(.a(new_n9716), .b(new_n9714), .O(new_n9717));
  inv1 g09524(.a(new_n9717), .O(\asquared[58] ));
  nor2 g09525(.a(new_n9704), .b(new_n9699), .O(new_n9719));
  nor2 g09526(.a(new_n9640), .b(new_n9447), .O(new_n9720));
  inv1 g09527(.a(new_n9720), .O(new_n9721));
  nor2 g09528(.a(new_n9442), .b(new_n9399), .O(new_n9722));
  inv1 g09529(.a(new_n9722), .O(new_n9723));
  nor2 g09530(.a(new_n9627), .b(new_n9576), .O(new_n9724));
  nor2 g09531(.a(new_n9570), .b(new_n9564), .O(new_n9725));
  inv1 g09532(.a(new_n9725), .O(new_n9726));
  nor2 g09533(.a(new_n9429), .b(new_n9423), .O(new_n9727));
  inv1 g09534(.a(new_n9727), .O(new_n9728));
  nor2 g09535(.a(new_n9728), .b(new_n9726), .O(new_n9729));
  nor2 g09536(.a(new_n9727), .b(new_n9725), .O(new_n9730));
  nor2 g09537(.a(new_n9730), .b(new_n9729), .O(new_n9731));
  nor2 g09538(.a(new_n9415), .b(new_n9409), .O(new_n9732));
  inv1 g09539(.a(new_n9732), .O(new_n9733));
  nor2 g09540(.a(new_n9733), .b(new_n9731), .O(new_n9734));
  inv1 g09541(.a(new_n9731), .O(new_n9735));
  nor2 g09542(.a(new_n9732), .b(new_n9735), .O(new_n9736));
  nor2 g09543(.a(new_n9736), .b(new_n9734), .O(new_n9737));
  inv1 g09544(.a(new_n9737), .O(new_n9738));
  nor2 g09545(.a(new_n9437), .b(new_n9432), .O(new_n9739));
  nor2 g09546(.a(new_n9739), .b(new_n9738), .O(new_n9740));
  inv1 g09547(.a(new_n9739), .O(new_n9741));
  nor2 g09548(.a(new_n9741), .b(new_n9737), .O(new_n9742));
  nor2 g09549(.a(new_n9742), .b(new_n9740), .O(new_n9743));
  inv1 g09550(.a(new_n9743), .O(new_n9744));
  nor2 g09551(.a(new_n9744), .b(new_n9724), .O(new_n9745));
  inv1 g09552(.a(new_n9724), .O(new_n9746));
  nor2 g09553(.a(new_n9743), .b(new_n9746), .O(new_n9747));
  nor2 g09554(.a(new_n9747), .b(new_n9745), .O(new_n9748));
  nor2 g09555(.a(new_n9748), .b(new_n9723), .O(new_n9749));
  inv1 g09556(.a(new_n9748), .O(new_n9750));
  nor2 g09557(.a(new_n9750), .b(new_n9722), .O(new_n9751));
  nor2 g09558(.a(new_n9751), .b(new_n9749), .O(new_n9752));
  inv1 g09559(.a(new_n9752), .O(new_n9753));
  nor2 g09560(.a(new_n9636), .b(new_n9631), .O(new_n9754));
  nor2 g09561(.a(new_n9754), .b(new_n9753), .O(new_n9755));
  inv1 g09562(.a(new_n9754), .O(new_n9756));
  nor2 g09563(.a(new_n9756), .b(new_n9752), .O(new_n9757));
  nor2 g09564(.a(new_n9757), .b(new_n9755), .O(new_n9758));
  nor2 g09565(.a(new_n9758), .b(new_n9721), .O(new_n9759));
  inv1 g09566(.a(new_n9758), .O(new_n9760));
  nor2 g09567(.a(new_n9760), .b(new_n9720), .O(new_n9761));
  nor2 g09568(.a(new_n9761), .b(new_n9759), .O(new_n9762));
  nor2 g09569(.a(new_n9694), .b(new_n9689), .O(new_n9763));
  inv1 g09570(.a(new_n9763), .O(new_n9764));
  nor2 g09571(.a(new_n9553), .b(new_n9550), .O(new_n9765));
  nor2 g09572(.a(new_n9658), .b(new_n194), .O(new_n9766));
  nor2 g09573(.a(new_n9766), .b(new_n9530), .O(new_n9767));
  inv1 g09574(.a(new_n9766), .O(new_n9768));
  nor2 g09575(.a(new_n9768), .b(new_n9531), .O(new_n9769));
  nor2 g09576(.a(new_n9769), .b(new_n9767), .O(new_n9770));
  nor2 g09577(.a(new_n9770), .b(new_n9667), .O(new_n9771));
  inv1 g09578(.a(new_n9667), .O(new_n9772));
  inv1 g09579(.a(new_n9770), .O(new_n9773));
  nor2 g09580(.a(new_n9773), .b(new_n9772), .O(new_n9774));
  nor2 g09581(.a(new_n9774), .b(new_n9771), .O(new_n9775));
  inv1 g09582(.a(new_n9775), .O(new_n9776));
  nor2 g09583(.a(new_n9536), .b(new_n9529), .O(new_n9777));
  inv1 g09584(.a(new_n9777), .O(new_n9778));
  nor2 g09585(.a(new_n9778), .b(new_n9776), .O(new_n9779));
  nor2 g09586(.a(new_n9777), .b(new_n9775), .O(new_n9780));
  nor2 g09587(.a(new_n9780), .b(new_n9779), .O(new_n9781));
  inv1 g09588(.a(new_n9781), .O(new_n9782));
  nor2 g09589(.a(new_n9498), .b(new_n9491), .O(new_n9783));
  nor2 g09590(.a(new_n9783), .b(new_n9782), .O(new_n9784));
  inv1 g09591(.a(new_n9783), .O(new_n9785));
  nor2 g09592(.a(new_n9785), .b(new_n9781), .O(new_n9786));
  nor2 g09593(.a(new_n9786), .b(new_n9784), .O(new_n9787));
  inv1 g09594(.a(new_n9787), .O(new_n9788));
  nor2 g09595(.a(new_n9545), .b(new_n9538), .O(new_n9789));
  nor2 g09596(.a(new_n9789), .b(new_n9788), .O(new_n9790));
  inv1 g09597(.a(new_n9789), .O(new_n9791));
  nor2 g09598(.a(new_n9791), .b(new_n9787), .O(new_n9792));
  nor2 g09599(.a(new_n9792), .b(new_n9790), .O(new_n9793));
  inv1 g09600(.a(new_n9793), .O(new_n9794));
  nor2 g09601(.a(new_n9794), .b(new_n9765), .O(new_n9795));
  inv1 g09602(.a(new_n9765), .O(new_n9796));
  nor2 g09603(.a(new_n9793), .b(new_n9796), .O(new_n9797));
  nor2 g09604(.a(new_n9797), .b(new_n9795), .O(new_n9798));
  inv1 g09605(.a(new_n9798), .O(new_n9799));
  nor2 g09606(.a(new_n9462), .b(new_n9455), .O(new_n9800));
  nor2 g09607(.a(new_n9589), .b(new_n9582), .O(new_n9801));
  nor2 g09608(.a(new_n9801), .b(new_n9800), .O(new_n9802));
  inv1 g09609(.a(new_n9800), .O(new_n9803));
  inv1 g09610(.a(new_n9801), .O(new_n9804));
  nor2 g09611(.a(new_n9804), .b(new_n9803), .O(new_n9805));
  nor2 g09612(.a(new_n9805), .b(new_n9802), .O(new_n9806));
  nor2 g09613(.a(new_n9615), .b(new_n9608), .O(new_n9807));
  nor2 g09614(.a(new_n9807), .b(new_n9806), .O(new_n9808));
  inv1 g09615(.a(new_n9806), .O(new_n9809));
  inv1 g09616(.a(new_n9807), .O(new_n9810));
  nor2 g09617(.a(new_n9810), .b(new_n9809), .O(new_n9811));
  nor2 g09618(.a(new_n9811), .b(new_n9808), .O(new_n9812));
  inv1 g09619(.a(new_n9812), .O(new_n9813));
  nor2 g09620(.a(new_n9489), .b(new_n9482), .O(new_n9814));
  nor2 g09621(.a(new_n9474), .b(new_n9467), .O(new_n9815));
  nor2 g09622(.a(new_n9815), .b(new_n9814), .O(new_n9816));
  inv1 g09623(.a(new_n9814), .O(new_n9817));
  inv1 g09624(.a(new_n9815), .O(new_n9818));
  nor2 g09625(.a(new_n9818), .b(new_n9817), .O(new_n9819));
  nor2 g09626(.a(new_n9819), .b(new_n9816), .O(new_n9820));
  nor2 g09627(.a(new_n9522), .b(new_n9515), .O(new_n9821));
  nor2 g09628(.a(new_n9821), .b(new_n9820), .O(new_n9822));
  inv1 g09629(.a(new_n9820), .O(new_n9823));
  inv1 g09630(.a(new_n9821), .O(new_n9824));
  nor2 g09631(.a(new_n9824), .b(new_n9823), .O(new_n9825));
  nor2 g09632(.a(new_n9825), .b(new_n9822), .O(new_n9826));
  inv1 g09633(.a(new_n9826), .O(new_n9827));
  nor2 g09634(.a(new_n9827), .b(new_n9813), .O(new_n9828));
  nor2 g09635(.a(new_n9826), .b(new_n9812), .O(new_n9829));
  nor2 g09636(.a(new_n9829), .b(new_n9828), .O(new_n9830));
  inv1 g09637(.a(new_n9830), .O(new_n9831));
  nor2 g09638(.a(new_n9624), .b(new_n9617), .O(new_n9832));
  nor2 g09639(.a(new_n9832), .b(new_n9831), .O(new_n9833));
  inv1 g09640(.a(new_n9832), .O(new_n9834));
  nor2 g09641(.a(new_n9834), .b(new_n9830), .O(new_n9835));
  nor2 g09642(.a(new_n9835), .b(new_n9833), .O(new_n9836));
  inv1 g09643(.a(new_n9836), .O(new_n9837));
  nor2 g09644(.a(new_n9837), .b(new_n9799), .O(new_n9838));
  nor2 g09645(.a(new_n9836), .b(new_n9798), .O(new_n9839));
  nor2 g09646(.a(new_n9839), .b(new_n9838), .O(new_n9840));
  nor2 g09647(.a(new_n9840), .b(new_n9764), .O(new_n9841));
  inv1 g09648(.a(new_n9840), .O(new_n9842));
  nor2 g09649(.a(new_n9842), .b(new_n9763), .O(new_n9843));
  nor2 g09650(.a(new_n9843), .b(new_n9841), .O(new_n9844));
  inv1 g09651(.a(new_n9844), .O(new_n9845));
  nor2 g09652(.a(new_n9395), .b(new_n9389), .O(new_n9846));
  inv1 g09653(.a(new_n9846), .O(new_n9847));
  nor2 g09654(.a(new_n4954), .b(new_n941), .O(new_n9848));
  inv1 g09655(.a(new_n9848), .O(new_n9849));
  nor2 g09656(.a(new_n6958), .b(new_n363), .O(new_n9850));
  nor2 g09657(.a(new_n5178), .b(new_n847), .O(new_n9851));
  nor2 g09658(.a(new_n9851), .b(new_n9850), .O(new_n9852));
  nor2 g09659(.a(new_n9597), .b(new_n7637), .O(new_n9853));
  nor2 g09660(.a(new_n9853), .b(new_n9852), .O(new_n9854));
  nor2 g09661(.a(new_n9854), .b(new_n9849), .O(new_n9855));
  inv1 g09662(.a(new_n9854), .O(new_n9856));
  nor2 g09663(.a(new_n9856), .b(new_n9848), .O(new_n9857));
  nor2 g09664(.a(new_n9857), .b(new_n9855), .O(new_n9858));
  inv1 g09665(.a(new_n9858), .O(new_n9859));
  nor2 g09666(.a(new_n8170), .b(new_n229), .O(new_n9860));
  inv1 g09667(.a(new_n9860), .O(new_n9861));
  nor2 g09668(.a(new_n4093), .b(new_n1425), .O(new_n9862));
  nor2 g09669(.a(new_n9862), .b(new_n9483), .O(new_n9863));
  inv1 g09670(.a(new_n9481), .O(new_n9864));
  nor2 g09671(.a(new_n4366), .b(new_n1425), .O(new_n9865));
  inv1 g09672(.a(new_n9865), .O(new_n9866));
  nor2 g09673(.a(new_n9866), .b(new_n9864), .O(new_n9867));
  nor2 g09674(.a(new_n9867), .b(new_n9863), .O(new_n9868));
  nor2 g09675(.a(new_n9868), .b(new_n9861), .O(new_n9869));
  inv1 g09676(.a(new_n9868), .O(new_n9870));
  nor2 g09677(.a(new_n9870), .b(new_n9860), .O(new_n9871));
  nor2 g09678(.a(new_n9871), .b(new_n9869), .O(new_n9872));
  inv1 g09679(.a(\a[58] ), .O(new_n9873));
  nor2 g09680(.a(new_n9873), .b(new_n198), .O(new_n9874));
  nor2 g09681(.a(new_n8476), .b(new_n214), .O(new_n9875));
  nor2 g09682(.a(new_n9875), .b(new_n9874), .O(new_n9876));
  inv1 g09683(.a(new_n9874), .O(new_n9877));
  inv1 g09684(.a(new_n9875), .O(new_n9878));
  nor2 g09685(.a(new_n9878), .b(new_n9877), .O(new_n9879));
  nor2 g09686(.a(new_n9879), .b(new_n9876), .O(new_n9880));
  nor2 g09687(.a(new_n9880), .b(new_n9161), .O(new_n9881));
  inv1 g09688(.a(new_n9880), .O(new_n9882));
  nor2 g09689(.a(new_n9882), .b(new_n9160), .O(new_n9883));
  nor2 g09690(.a(new_n9883), .b(new_n9881), .O(new_n9884));
  nor2 g09691(.a(new_n9884), .b(new_n9872), .O(new_n9885));
  inv1 g09692(.a(new_n9872), .O(new_n9886));
  inv1 g09693(.a(new_n9884), .O(new_n9887));
  nor2 g09694(.a(new_n9887), .b(new_n9886), .O(new_n9888));
  nor2 g09695(.a(new_n9888), .b(new_n9885), .O(new_n9889));
  nor2 g09696(.a(new_n9889), .b(new_n9859), .O(new_n9890));
  inv1 g09697(.a(new_n9889), .O(new_n9891));
  nor2 g09698(.a(new_n9891), .b(new_n9858), .O(new_n9892));
  nor2 g09699(.a(new_n9892), .b(new_n9890), .O(new_n9893));
  inv1 g09700(.a(new_n9893), .O(new_n9894));
  nor2 g09701(.a(new_n3231), .b(new_n1903), .O(new_n9895));
  inv1 g09702(.a(new_n9895), .O(new_n9896));
  nor2 g09703(.a(new_n2826), .b(new_n2184), .O(new_n9897));
  nor2 g09704(.a(new_n9897), .b(new_n9583), .O(new_n9898));
  nor2 g09705(.a(new_n3057), .b(new_n2184), .O(new_n9899));
  inv1 g09706(.a(new_n9899), .O(new_n9900));
  nor2 g09707(.a(new_n9900), .b(new_n9135), .O(new_n9901));
  nor2 g09708(.a(new_n9901), .b(new_n9898), .O(new_n9902));
  nor2 g09709(.a(new_n9902), .b(new_n9896), .O(new_n9903));
  inv1 g09710(.a(new_n9902), .O(new_n9904));
  nor2 g09711(.a(new_n9904), .b(new_n9895), .O(new_n9905));
  nor2 g09712(.a(new_n9905), .b(new_n9903), .O(new_n9906));
  inv1 g09713(.a(new_n9906), .O(new_n9907));
  nor2 g09714(.a(new_n4682), .b(new_n1086), .O(new_n9908));
  nor2 g09715(.a(new_n7537), .b(new_n295), .O(new_n9909));
  nor2 g09716(.a(new_n7294), .b(new_n322), .O(new_n9910));
  nor2 g09717(.a(new_n9910), .b(new_n9909), .O(new_n9911));
  nor2 g09718(.a(new_n7537), .b(new_n322), .O(new_n9912));
  inv1 g09719(.a(new_n9912), .O(new_n9913));
  nor2 g09720(.a(new_n9913), .b(new_n9602), .O(new_n9914));
  nor2 g09721(.a(new_n9914), .b(new_n9911), .O(new_n9915));
  inv1 g09722(.a(new_n9915), .O(new_n9916));
  nor2 g09723(.a(new_n9916), .b(new_n9908), .O(new_n9917));
  inv1 g09724(.a(new_n9908), .O(new_n9918));
  nor2 g09725(.a(new_n9915), .b(new_n9918), .O(new_n9919));
  nor2 g09726(.a(new_n9919), .b(new_n9917), .O(new_n9920));
  nor2 g09727(.a(new_n3870), .b(new_n1493), .O(new_n9921));
  inv1 g09728(.a(new_n9921), .O(new_n9922));
  nor2 g09729(.a(new_n3533), .b(new_n1736), .O(new_n9923));
  nor2 g09730(.a(new_n9923), .b(new_n9609), .O(new_n9924));
  nor2 g09731(.a(new_n3722), .b(new_n1736), .O(new_n9925));
  inv1 g09732(.a(new_n9925), .O(new_n9926));
  nor2 g09733(.a(new_n9926), .b(new_n9122), .O(new_n9927));
  nor2 g09734(.a(new_n9927), .b(new_n9924), .O(new_n9928));
  nor2 g09735(.a(new_n9928), .b(new_n9922), .O(new_n9929));
  inv1 g09736(.a(new_n9928), .O(new_n9930));
  nor2 g09737(.a(new_n9930), .b(new_n9921), .O(new_n9931));
  nor2 g09738(.a(new_n9931), .b(new_n9929), .O(new_n9932));
  nor2 g09739(.a(new_n9932), .b(new_n9920), .O(new_n9933));
  inv1 g09740(.a(new_n9920), .O(new_n9934));
  inv1 g09741(.a(new_n9932), .O(new_n9935));
  nor2 g09742(.a(new_n9935), .b(new_n9934), .O(new_n9936));
  nor2 g09743(.a(new_n9936), .b(new_n9933), .O(new_n9937));
  nor2 g09744(.a(new_n9937), .b(new_n9907), .O(new_n9938));
  inv1 g09745(.a(new_n9937), .O(new_n9939));
  nor2 g09746(.a(new_n9939), .b(new_n9906), .O(new_n9940));
  nor2 g09747(.a(new_n9940), .b(new_n9938), .O(new_n9941));
  inv1 g09748(.a(new_n9941), .O(new_n9942));
  nor2 g09749(.a(new_n9942), .b(new_n9894), .O(new_n9943));
  nor2 g09750(.a(new_n9941), .b(new_n9893), .O(new_n9944));
  nor2 g09751(.a(new_n9944), .b(new_n9943), .O(new_n9945));
  nor2 g09752(.a(new_n9945), .b(new_n9847), .O(new_n9946));
  inv1 g09753(.a(new_n9945), .O(new_n9947));
  nor2 g09754(.a(new_n9947), .b(new_n9846), .O(new_n9948));
  nor2 g09755(.a(new_n9948), .b(new_n9946), .O(new_n9949));
  inv1 g09756(.a(new_n9949), .O(new_n9950));
  nor2 g09757(.a(new_n9685), .b(new_n9652), .O(new_n9951));
  nor2 g09758(.a(new_n9511), .b(new_n9504), .O(new_n9952));
  nor2 g09759(.a(new_n9601), .b(new_n9595), .O(new_n9953));
  nor2 g09760(.a(new_n9953), .b(new_n9952), .O(new_n9954));
  inv1 g09761(.a(new_n9952), .O(new_n9955));
  inv1 g09762(.a(new_n9953), .O(new_n9956));
  nor2 g09763(.a(new_n9956), .b(new_n9955), .O(new_n9957));
  nor2 g09764(.a(new_n9957), .b(new_n9954), .O(new_n9958));
  nor2 g09765(.a(new_n9671), .b(new_n9661), .O(new_n9959));
  inv1 g09766(.a(new_n9959), .O(new_n9960));
  nor2 g09767(.a(new_n9960), .b(new_n9958), .O(new_n9961));
  inv1 g09768(.a(new_n9958), .O(new_n9962));
  nor2 g09769(.a(new_n9959), .b(new_n9962), .O(new_n9963));
  nor2 g09770(.a(new_n9963), .b(new_n9961), .O(new_n9964));
  nor2 g09771(.a(new_n9682), .b(new_n9676), .O(new_n9965));
  inv1 g09772(.a(new_n9965), .O(new_n9966));
  nor2 g09773(.a(new_n9966), .b(new_n9964), .O(new_n9967));
  inv1 g09774(.a(new_n9964), .O(new_n9968));
  nor2 g09775(.a(new_n9965), .b(new_n9968), .O(new_n9969));
  nor2 g09776(.a(new_n9969), .b(new_n9967), .O(new_n9970));
  nor2 g09777(.a(new_n8946), .b(new_n203), .O(new_n9971));
  inv1 g09778(.a(new_n9971), .O(new_n9972));
  nor2 g09779(.a(new_n4425), .b(new_n1199), .O(new_n9973));
  nor2 g09780(.a(new_n8026), .b(new_n257), .O(new_n9974));
  nor2 g09781(.a(new_n9974), .b(new_n9973), .O(new_n9975));
  inv1 g09782(.a(new_n9973), .O(new_n9976));
  inv1 g09783(.a(new_n9974), .O(new_n9977));
  nor2 g09784(.a(new_n9977), .b(new_n9976), .O(new_n9978));
  nor2 g09785(.a(new_n9978), .b(new_n9975), .O(new_n9979));
  nor2 g09786(.a(new_n9979), .b(new_n9972), .O(new_n9980));
  inv1 g09787(.a(new_n9979), .O(new_n9981));
  nor2 g09788(.a(new_n9981), .b(new_n9971), .O(new_n9982));
  nor2 g09789(.a(new_n9982), .b(new_n9980), .O(new_n9983));
  inv1 g09790(.a(new_n9983), .O(new_n9984));
  nor2 g09791(.a(new_n6570), .b(new_n502), .O(new_n9985));
  nor2 g09792(.a(new_n9985), .b(new_n6492), .O(new_n9986));
  inv1 g09793(.a(new_n8593), .O(new_n9987));
  nor2 g09794(.a(new_n6570), .b(new_n800), .O(new_n9988));
  inv1 g09795(.a(new_n9988), .O(new_n9989));
  nor2 g09796(.a(new_n9989), .b(new_n9987), .O(new_n9990));
  nor2 g09797(.a(new_n9990), .b(new_n9986), .O(new_n9991));
  inv1 g09798(.a(new_n9991), .O(new_n9992));
  nor2 g09799(.a(new_n9992), .b(new_n9456), .O(new_n9993));
  nor2 g09800(.a(new_n9991), .b(new_n9457), .O(new_n9994));
  nor2 g09801(.a(new_n9994), .b(new_n9993), .O(new_n9995));
  nor2 g09802(.a(new_n5971), .b(new_n613), .O(new_n9996));
  nor2 g09803(.a(new_n6274), .b(new_n569), .O(new_n9997));
  nor2 g09804(.a(new_n9997), .b(new_n9996), .O(new_n9998));
  nor2 g09805(.a(new_n9526), .b(new_n9518), .O(new_n9999));
  nor2 g09806(.a(new_n9999), .b(new_n9998), .O(new_n10000));
  nor2 g09807(.a(new_n10000), .b(new_n8201), .O(new_n10001));
  inv1 g09808(.a(new_n10000), .O(new_n10002));
  nor2 g09809(.a(new_n10002), .b(new_n8200), .O(new_n10003));
  nor2 g09810(.a(new_n10003), .b(new_n10001), .O(new_n10004));
  nor2 g09811(.a(new_n10004), .b(new_n9995), .O(new_n10005));
  inv1 g09812(.a(new_n9995), .O(new_n10006));
  inv1 g09813(.a(new_n10004), .O(new_n10007));
  nor2 g09814(.a(new_n10007), .b(new_n10006), .O(new_n10008));
  nor2 g09815(.a(new_n10008), .b(new_n10005), .O(new_n10009));
  nor2 g09816(.a(new_n10009), .b(new_n9984), .O(new_n10010));
  inv1 g09817(.a(new_n10009), .O(new_n10011));
  nor2 g09818(.a(new_n10011), .b(new_n9983), .O(new_n10012));
  nor2 g09819(.a(new_n10012), .b(new_n10010), .O(new_n10013));
  nor2 g09820(.a(new_n10013), .b(new_n9970), .O(new_n10014));
  inv1 g09821(.a(new_n9970), .O(new_n10015));
  inv1 g09822(.a(new_n10013), .O(new_n10016));
  nor2 g09823(.a(new_n10016), .b(new_n10015), .O(new_n10017));
  nor2 g09824(.a(new_n10017), .b(new_n10014), .O(new_n10018));
  inv1 g09825(.a(new_n10018), .O(new_n10019));
  nor2 g09826(.a(new_n10019), .b(new_n9951), .O(new_n10020));
  inv1 g09827(.a(new_n9951), .O(new_n10021));
  nor2 g09828(.a(new_n10018), .b(new_n10021), .O(new_n10022));
  nor2 g09829(.a(new_n10022), .b(new_n10020), .O(new_n10023));
  inv1 g09830(.a(new_n10023), .O(new_n10024));
  nor2 g09831(.a(new_n10024), .b(new_n9950), .O(new_n10025));
  nor2 g09832(.a(new_n10023), .b(new_n9949), .O(new_n10026));
  nor2 g09833(.a(new_n10026), .b(new_n10025), .O(new_n10027));
  inv1 g09834(.a(new_n10027), .O(new_n10028));
  nor2 g09835(.a(new_n10028), .b(new_n9845), .O(new_n10029));
  nor2 g09836(.a(new_n10027), .b(new_n9844), .O(new_n10030));
  nor2 g09837(.a(new_n10030), .b(new_n10029), .O(new_n10031));
  nor2 g09838(.a(new_n10031), .b(new_n9762), .O(new_n10032));
  inv1 g09839(.a(new_n9762), .O(new_n10033));
  inv1 g09840(.a(new_n10031), .O(new_n10034));
  nor2 g09841(.a(new_n10034), .b(new_n10033), .O(new_n10035));
  nor2 g09842(.a(new_n10035), .b(new_n10032), .O(new_n10036));
  inv1 g09843(.a(new_n10036), .O(new_n10037));
  nor2 g09844(.a(new_n10037), .b(new_n9719), .O(new_n10038));
  inv1 g09845(.a(new_n9719), .O(new_n10039));
  nor2 g09846(.a(new_n10036), .b(new_n10039), .O(new_n10040));
  nor2 g09847(.a(new_n10040), .b(new_n10038), .O(new_n10041));
  inv1 g09848(.a(new_n10041), .O(new_n10042));
  nor2 g09849(.a(new_n9714), .b(new_n9710), .O(new_n10043));
  nor2 g09850(.a(new_n10043), .b(new_n10042), .O(new_n10044));
  inv1 g09851(.a(new_n10043), .O(new_n10045));
  nor2 g09852(.a(new_n10045), .b(new_n10041), .O(new_n10046));
  nor2 g09853(.a(new_n10046), .b(new_n10044), .O(new_n10047));
  inv1 g09854(.a(new_n10047), .O(\asquared[59] ));
  nor2 g09855(.a(new_n10029), .b(new_n9843), .O(new_n10049));
  inv1 g09856(.a(new_n10049), .O(new_n10050));
  nor2 g09857(.a(new_n10025), .b(new_n10020), .O(new_n10051));
  nor2 g09858(.a(new_n9838), .b(new_n9795), .O(new_n10052));
  nor2 g09859(.a(new_n10017), .b(new_n9969), .O(new_n10053));
  nor2 g09860(.a(new_n9963), .b(new_n9957), .O(new_n10054));
  inv1 g09861(.a(new_n10054), .O(new_n10055));
  nor2 g09862(.a(new_n9825), .b(new_n9819), .O(new_n10056));
  inv1 g09863(.a(new_n10056), .O(new_n10057));
  nor2 g09864(.a(new_n10057), .b(new_n10055), .O(new_n10058));
  nor2 g09865(.a(new_n10056), .b(new_n10054), .O(new_n10059));
  nor2 g09866(.a(new_n10059), .b(new_n10058), .O(new_n10060));
  nor2 g09867(.a(new_n9811), .b(new_n9805), .O(new_n10061));
  inv1 g09868(.a(new_n10061), .O(new_n10062));
  nor2 g09869(.a(new_n10062), .b(new_n10060), .O(new_n10063));
  inv1 g09870(.a(new_n10060), .O(new_n10064));
  nor2 g09871(.a(new_n10061), .b(new_n10064), .O(new_n10065));
  nor2 g09872(.a(new_n10065), .b(new_n10063), .O(new_n10066));
  inv1 g09873(.a(new_n10066), .O(new_n10067));
  nor2 g09874(.a(new_n9833), .b(new_n9828), .O(new_n10068));
  nor2 g09875(.a(new_n10068), .b(new_n10067), .O(new_n10069));
  inv1 g09876(.a(new_n10068), .O(new_n10070));
  nor2 g09877(.a(new_n10070), .b(new_n10066), .O(new_n10071));
  nor2 g09878(.a(new_n10071), .b(new_n10069), .O(new_n10072));
  inv1 g09879(.a(new_n10072), .O(new_n10073));
  nor2 g09880(.a(new_n10073), .b(new_n10053), .O(new_n10074));
  inv1 g09881(.a(new_n10053), .O(new_n10075));
  nor2 g09882(.a(new_n10072), .b(new_n10075), .O(new_n10076));
  nor2 g09883(.a(new_n10076), .b(new_n10074), .O(new_n10077));
  inv1 g09884(.a(new_n10077), .O(new_n10078));
  nor2 g09885(.a(new_n10078), .b(new_n10052), .O(new_n10079));
  inv1 g09886(.a(new_n10052), .O(new_n10080));
  nor2 g09887(.a(new_n10077), .b(new_n10080), .O(new_n10081));
  nor2 g09888(.a(new_n10081), .b(new_n10079), .O(new_n10082));
  inv1 g09889(.a(new_n10082), .O(new_n10083));
  nor2 g09890(.a(new_n10083), .b(new_n10051), .O(new_n10084));
  inv1 g09891(.a(new_n10051), .O(new_n10085));
  nor2 g09892(.a(new_n10082), .b(new_n10085), .O(new_n10086));
  nor2 g09893(.a(new_n10086), .b(new_n10084), .O(new_n10087));
  nor2 g09894(.a(new_n10087), .b(new_n10050), .O(new_n10088));
  inv1 g09895(.a(new_n10087), .O(new_n10089));
  nor2 g09896(.a(new_n10089), .b(new_n10049), .O(new_n10090));
  nor2 g09897(.a(new_n10090), .b(new_n10088), .O(new_n10091));
  inv1 g09898(.a(new_n10091), .O(new_n10092));
  nor2 g09899(.a(new_n9755), .b(new_n9751), .O(new_n10093));
  nor2 g09900(.a(new_n9940), .b(new_n9933), .O(new_n10094));
  inv1 g09901(.a(new_n10094), .O(new_n10095));
  nor2 g09902(.a(new_n10012), .b(new_n10005), .O(new_n10096));
  inv1 g09903(.a(new_n10096), .O(new_n10097));
  nor2 g09904(.a(new_n10097), .b(new_n10095), .O(new_n10098));
  nor2 g09905(.a(new_n10096), .b(new_n10094), .O(new_n10099));
  nor2 g09906(.a(new_n10099), .b(new_n10098), .O(new_n10100));
  nor2 g09907(.a(new_n9892), .b(new_n9885), .O(new_n10101));
  inv1 g09908(.a(new_n10101), .O(new_n10102));
  nor2 g09909(.a(new_n10102), .b(new_n10100), .O(new_n10103));
  inv1 g09910(.a(new_n10100), .O(new_n10104));
  nor2 g09911(.a(new_n10101), .b(new_n10104), .O(new_n10105));
  nor2 g09912(.a(new_n10105), .b(new_n10103), .O(new_n10106));
  inv1 g09913(.a(new_n10106), .O(new_n10107));
  nor2 g09914(.a(new_n9948), .b(new_n9943), .O(new_n10108));
  nor2 g09915(.a(new_n9883), .b(new_n9876), .O(new_n10109));
  nor2 g09916(.a(new_n9982), .b(new_n9975), .O(new_n10110));
  nor2 g09917(.a(new_n10110), .b(new_n10109), .O(new_n10111));
  inv1 g09918(.a(new_n10109), .O(new_n10112));
  inv1 g09919(.a(new_n10110), .O(new_n10113));
  nor2 g09920(.a(new_n10113), .b(new_n10112), .O(new_n10114));
  nor2 g09921(.a(new_n10114), .b(new_n10111), .O(new_n10115));
  nor2 g09922(.a(new_n9857), .b(new_n9852), .O(new_n10116));
  nor2 g09923(.a(new_n10116), .b(new_n10115), .O(new_n10117));
  inv1 g09924(.a(new_n10115), .O(new_n10118));
  inv1 g09925(.a(new_n10116), .O(new_n10119));
  nor2 g09926(.a(new_n10119), .b(new_n10118), .O(new_n10120));
  nor2 g09927(.a(new_n10120), .b(new_n10117), .O(new_n10121));
  inv1 g09928(.a(new_n10121), .O(new_n10122));
  nor2 g09929(.a(new_n9871), .b(new_n9863), .O(new_n10123));
  nor2 g09930(.a(new_n9931), .b(new_n9924), .O(new_n10124));
  nor2 g09931(.a(new_n10124), .b(new_n10123), .O(new_n10125));
  inv1 g09932(.a(new_n10123), .O(new_n10126));
  inv1 g09933(.a(new_n10124), .O(new_n10127));
  nor2 g09934(.a(new_n10127), .b(new_n10126), .O(new_n10128));
  nor2 g09935(.a(new_n10128), .b(new_n10125), .O(new_n10129));
  nor2 g09936(.a(new_n9917), .b(new_n9911), .O(new_n10130));
  nor2 g09937(.a(new_n10130), .b(new_n10129), .O(new_n10131));
  inv1 g09938(.a(new_n10129), .O(new_n10132));
  inv1 g09939(.a(new_n10130), .O(new_n10133));
  nor2 g09940(.a(new_n10133), .b(new_n10132), .O(new_n10134));
  nor2 g09941(.a(new_n10134), .b(new_n10131), .O(new_n10135));
  inv1 g09942(.a(new_n10135), .O(new_n10136));
  nor2 g09943(.a(new_n2937), .b(new_n9873), .O(new_n10137));
  nor2 g09944(.a(new_n9873), .b(new_n194), .O(new_n10138));
  nor2 g09945(.a(new_n10138), .b(\a[30] ), .O(new_n10139));
  nor2 g09946(.a(new_n10139), .b(new_n10137), .O(new_n10140));
  nor2 g09947(.a(new_n10003), .b(new_n9998), .O(new_n10141));
  nor2 g09948(.a(new_n10141), .b(new_n10140), .O(new_n10142));
  inv1 g09949(.a(new_n10140), .O(new_n10143));
  inv1 g09950(.a(new_n10141), .O(new_n10144));
  nor2 g09951(.a(new_n10144), .b(new_n10143), .O(new_n10145));
  nor2 g09952(.a(new_n10145), .b(new_n10142), .O(new_n10146));
  inv1 g09953(.a(new_n10146), .O(new_n10147));
  nor2 g09954(.a(new_n9993), .b(new_n9986), .O(new_n10148));
  inv1 g09955(.a(new_n10148), .O(new_n10149));
  nor2 g09956(.a(new_n10149), .b(new_n10147), .O(new_n10150));
  nor2 g09957(.a(new_n10148), .b(new_n10146), .O(new_n10151));
  nor2 g09958(.a(new_n10151), .b(new_n10150), .O(new_n10152));
  inv1 g09959(.a(new_n10152), .O(new_n10153));
  nor2 g09960(.a(new_n10153), .b(new_n10136), .O(new_n10154));
  nor2 g09961(.a(new_n10152), .b(new_n10135), .O(new_n10155));
  nor2 g09962(.a(new_n10155), .b(new_n10154), .O(new_n10156));
  inv1 g09963(.a(new_n10156), .O(new_n10157));
  nor2 g09964(.a(new_n10157), .b(new_n10122), .O(new_n10158));
  nor2 g09965(.a(new_n10156), .b(new_n10121), .O(new_n10159));
  nor2 g09966(.a(new_n10159), .b(new_n10158), .O(new_n10160));
  inv1 g09967(.a(new_n10160), .O(new_n10161));
  nor2 g09968(.a(new_n10161), .b(new_n10108), .O(new_n10162));
  inv1 g09969(.a(new_n10108), .O(new_n10163));
  nor2 g09970(.a(new_n10160), .b(new_n10163), .O(new_n10164));
  nor2 g09971(.a(new_n10164), .b(new_n10162), .O(new_n10165));
  inv1 g09972(.a(new_n10165), .O(new_n10166));
  nor2 g09973(.a(new_n10166), .b(new_n10107), .O(new_n10167));
  nor2 g09974(.a(new_n10165), .b(new_n10106), .O(new_n10168));
  nor2 g09975(.a(new_n10168), .b(new_n10167), .O(new_n10169));
  inv1 g09976(.a(new_n10169), .O(new_n10170));
  nor2 g09977(.a(new_n10170), .b(new_n10093), .O(new_n10171));
  inv1 g09978(.a(new_n10093), .O(new_n10172));
  nor2 g09979(.a(new_n10169), .b(new_n10172), .O(new_n10173));
  nor2 g09980(.a(new_n10173), .b(new_n10171), .O(new_n10174));
  inv1 g09981(.a(new_n10174), .O(new_n10175));
  nor2 g09982(.a(new_n9745), .b(new_n9740), .O(new_n10176));
  inv1 g09983(.a(new_n10176), .O(new_n10177));
  nor2 g09984(.a(new_n9790), .b(new_n9784), .O(new_n10178));
  nor2 g09985(.a(new_n8476), .b(new_n229), .O(new_n10179));
  nor2 g09986(.a(new_n4682), .b(new_n1199), .O(new_n10180));
  nor2 g09987(.a(new_n10180), .b(new_n10179), .O(new_n10181));
  inv1 g09988(.a(new_n10179), .O(new_n10182));
  inv1 g09989(.a(new_n10180), .O(new_n10183));
  nor2 g09990(.a(new_n10183), .b(new_n10182), .O(new_n10184));
  nor2 g09991(.a(new_n10184), .b(new_n10181), .O(new_n10185));
  nor2 g09992(.a(new_n10185), .b(new_n9470), .O(new_n10186));
  inv1 g09993(.a(new_n10185), .O(new_n10187));
  nor2 g09994(.a(new_n10187), .b(new_n9469), .O(new_n10188));
  nor2 g09995(.a(new_n10188), .b(new_n10186), .O(new_n10189));
  nor2 g09996(.a(new_n9658), .b(new_n196), .O(new_n10190));
  nor2 g09997(.a(new_n9156), .b(new_n203), .O(new_n10191));
  nor2 g09998(.a(new_n10191), .b(new_n10190), .O(new_n10192));
  nor2 g09999(.a(new_n9658), .b(new_n203), .O(new_n10193));
  inv1 g10000(.a(new_n10193), .O(new_n10194));
  nor2 g10001(.a(new_n10194), .b(new_n9161), .O(new_n10195));
  nor2 g10002(.a(new_n10195), .b(new_n10192), .O(new_n10196));
  inv1 g10003(.a(new_n10196), .O(new_n10197));
  nor2 g10004(.a(new_n10197), .b(new_n9769), .O(new_n10198));
  inv1 g10005(.a(new_n9769), .O(new_n10199));
  nor2 g10006(.a(new_n10196), .b(new_n10199), .O(new_n10200));
  nor2 g10007(.a(new_n10200), .b(new_n10198), .O(new_n10201));
  nor2 g10008(.a(new_n9905), .b(new_n9898), .O(new_n10202));
  inv1 g10009(.a(new_n10202), .O(new_n10203));
  nor2 g10010(.a(new_n10203), .b(new_n10201), .O(new_n10204));
  inv1 g10011(.a(new_n10201), .O(new_n10205));
  nor2 g10012(.a(new_n10202), .b(new_n10205), .O(new_n10206));
  nor2 g10013(.a(new_n10206), .b(new_n10204), .O(new_n10207));
  inv1 g10014(.a(new_n10207), .O(new_n10208));
  nor2 g10015(.a(new_n10208), .b(new_n10189), .O(new_n10209));
  inv1 g10016(.a(new_n10189), .O(new_n10210));
  nor2 g10017(.a(new_n10207), .b(new_n10210), .O(new_n10211));
  nor2 g10018(.a(new_n10211), .b(new_n10209), .O(new_n10212));
  nor2 g10019(.a(new_n5393), .b(new_n847), .O(new_n10213));
  nor2 g10020(.a(new_n5178), .b(new_n941), .O(new_n10214));
  nor2 g10021(.a(new_n10214), .b(new_n10213), .O(new_n10215));
  inv1 g10022(.a(new_n9851), .O(new_n10216));
  nor2 g10023(.a(new_n5393), .b(new_n941), .O(new_n10217));
  inv1 g10024(.a(new_n10217), .O(new_n10218));
  nor2 g10025(.a(new_n10218), .b(new_n10216), .O(new_n10219));
  nor2 g10026(.a(new_n10219), .b(new_n10215), .O(new_n10220));
  nor2 g10027(.a(new_n10220), .b(new_n9913), .O(new_n10221));
  inv1 g10028(.a(new_n10220), .O(new_n10222));
  nor2 g10029(.a(new_n10222), .b(new_n9912), .O(new_n10223));
  nor2 g10030(.a(new_n10223), .b(new_n10221), .O(new_n10224));
  inv1 g10031(.a(new_n10224), .O(new_n10225));
  nor2 g10032(.a(new_n6893), .b(new_n502), .O(new_n10226));
  nor2 g10033(.a(new_n6570), .b(new_n569), .O(new_n10227));
  nor2 g10034(.a(new_n10227), .b(new_n7598), .O(new_n10228));
  nor2 g10035(.a(new_n6570), .b(new_n699), .O(new_n10229));
  inv1 g10036(.a(new_n10229), .O(new_n10230));
  nor2 g10037(.a(new_n10230), .b(new_n9526), .O(new_n10231));
  nor2 g10038(.a(new_n10231), .b(new_n10228), .O(new_n10232));
  inv1 g10039(.a(new_n10232), .O(new_n10233));
  nor2 g10040(.a(new_n10233), .b(new_n10226), .O(new_n10234));
  inv1 g10041(.a(new_n10226), .O(new_n10235));
  nor2 g10042(.a(new_n10232), .b(new_n10235), .O(new_n10236));
  nor2 g10043(.a(new_n10236), .b(new_n10234), .O(new_n10237));
  nor2 g10044(.a(new_n2660), .b(new_n2506), .O(new_n10238));
  nor2 g10045(.a(new_n2826), .b(new_n2433), .O(new_n10239));
  nor2 g10046(.a(new_n10239), .b(new_n10238), .O(new_n10240));
  inv1 g10047(.a(new_n10238), .O(new_n10241));
  inv1 g10048(.a(new_n10239), .O(new_n10242));
  nor2 g10049(.a(new_n10242), .b(new_n10241), .O(new_n10243));
  nor2 g10050(.a(new_n10243), .b(new_n10240), .O(new_n10244));
  nor2 g10051(.a(new_n10244), .b(new_n9518), .O(new_n10245));
  inv1 g10052(.a(new_n10244), .O(new_n10246));
  nor2 g10053(.a(new_n10246), .b(new_n9517), .O(new_n10247));
  nor2 g10054(.a(new_n10247), .b(new_n10245), .O(new_n10248));
  nor2 g10055(.a(new_n10248), .b(new_n10237), .O(new_n10249));
  inv1 g10056(.a(new_n10237), .O(new_n10250));
  inv1 g10057(.a(new_n10248), .O(new_n10251));
  nor2 g10058(.a(new_n10251), .b(new_n10250), .O(new_n10252));
  nor2 g10059(.a(new_n10252), .b(new_n10249), .O(new_n10253));
  nor2 g10060(.a(new_n10253), .b(new_n10225), .O(new_n10254));
  inv1 g10061(.a(new_n10253), .O(new_n10255));
  nor2 g10062(.a(new_n10255), .b(new_n10224), .O(new_n10256));
  nor2 g10063(.a(new_n10256), .b(new_n10254), .O(new_n10257));
  nor2 g10064(.a(new_n10257), .b(new_n10212), .O(new_n10258));
  inv1 g10065(.a(new_n10212), .O(new_n10259));
  inv1 g10066(.a(new_n10257), .O(new_n10260));
  nor2 g10067(.a(new_n10260), .b(new_n10259), .O(new_n10261));
  nor2 g10068(.a(new_n10261), .b(new_n10258), .O(new_n10262));
  inv1 g10069(.a(new_n10262), .O(new_n10263));
  nor2 g10070(.a(new_n10263), .b(new_n10178), .O(new_n10264));
  inv1 g10071(.a(new_n10178), .O(new_n10265));
  nor2 g10072(.a(new_n10262), .b(new_n10265), .O(new_n10266));
  nor2 g10073(.a(new_n10266), .b(new_n10264), .O(new_n10267));
  nor2 g10074(.a(new_n10267), .b(new_n10177), .O(new_n10268));
  inv1 g10075(.a(new_n10267), .O(new_n10269));
  nor2 g10076(.a(new_n10269), .b(new_n10176), .O(new_n10270));
  nor2 g10077(.a(new_n10270), .b(new_n10268), .O(new_n10271));
  inv1 g10078(.a(new_n10271), .O(new_n10272));
  nor2 g10079(.a(new_n9779), .b(new_n9774), .O(new_n10273));
  inv1 g10080(.a(new_n10273), .O(new_n10274));
  nor2 g10081(.a(new_n8170), .b(new_n257), .O(new_n10275));
  nor2 g10082(.a(new_n8026), .b(new_n295), .O(new_n10276));
  nor2 g10083(.a(new_n4954), .b(new_n1086), .O(new_n10277));
  nor2 g10084(.a(new_n10277), .b(new_n10276), .O(new_n10278));
  nor2 g10085(.a(new_n8026), .b(new_n1086), .O(new_n10279));
  inv1 g10086(.a(new_n10279), .O(new_n10280));
  nor2 g10087(.a(new_n10280), .b(new_n6700), .O(new_n10281));
  nor2 g10088(.a(new_n10281), .b(new_n10278), .O(new_n10282));
  inv1 g10089(.a(new_n10282), .O(new_n10283));
  nor2 g10090(.a(new_n10283), .b(new_n10275), .O(new_n10284));
  inv1 g10091(.a(new_n10275), .O(new_n10285));
  nor2 g10092(.a(new_n10282), .b(new_n10285), .O(new_n10286));
  nor2 g10093(.a(new_n10286), .b(new_n10284), .O(new_n10287));
  nor2 g10094(.a(new_n7294), .b(new_n363), .O(new_n10288));
  inv1 g10095(.a(new_n10288), .O(new_n10289));
  nor2 g10096(.a(new_n5796), .b(new_n800), .O(new_n10290));
  nor2 g10097(.a(new_n6958), .b(new_n438), .O(new_n10291));
  nor2 g10098(.a(new_n10291), .b(new_n10290), .O(new_n10292));
  inv1 g10099(.a(new_n8659), .O(new_n10293));
  nor2 g10100(.a(new_n6958), .b(new_n800), .O(new_n10294));
  inv1 g10101(.a(new_n10294), .O(new_n10295));
  nor2 g10102(.a(new_n10295), .b(new_n10293), .O(new_n10296));
  nor2 g10103(.a(new_n10296), .b(new_n10292), .O(new_n10297));
  nor2 g10104(.a(new_n10297), .b(new_n10289), .O(new_n10298));
  inv1 g10105(.a(new_n10297), .O(new_n10299));
  nor2 g10106(.a(new_n10299), .b(new_n10288), .O(new_n10300));
  nor2 g10107(.a(new_n10300), .b(new_n10298), .O(new_n10301));
  nor2 g10108(.a(new_n10301), .b(new_n10287), .O(new_n10302));
  inv1 g10109(.a(new_n10287), .O(new_n10303));
  inv1 g10110(.a(new_n10301), .O(new_n10304));
  nor2 g10111(.a(new_n10304), .b(new_n10303), .O(new_n10305));
  nor2 g10112(.a(new_n10305), .b(new_n10302), .O(new_n10306));
  nor2 g10113(.a(new_n10306), .b(new_n10274), .O(new_n10307));
  inv1 g10114(.a(new_n10306), .O(new_n10308));
  nor2 g10115(.a(new_n10308), .b(new_n10273), .O(new_n10309));
  nor2 g10116(.a(new_n10309), .b(new_n10307), .O(new_n10310));
  nor2 g10117(.a(new_n9736), .b(new_n9730), .O(new_n10311));
  inv1 g10118(.a(new_n10311), .O(new_n10312));
  nor2 g10119(.a(new_n10312), .b(new_n10310), .O(new_n10313));
  inv1 g10120(.a(new_n10310), .O(new_n10314));
  nor2 g10121(.a(new_n10311), .b(new_n10314), .O(new_n10315));
  nor2 g10122(.a(new_n10315), .b(new_n10313), .O(new_n10316));
  inv1 g10123(.a(new_n10316), .O(new_n10317));
  nor2 g10124(.a(new_n3231), .b(new_n2121), .O(new_n10318));
  inv1 g10125(.a(new_n10318), .O(new_n10319));
  inv1 g10126(.a(\a[59] ), .O(new_n10320));
  nor2 g10127(.a(new_n10320), .b(new_n198), .O(new_n10321));
  nor2 g10128(.a(new_n10321), .b(new_n9899), .O(new_n10322));
  inv1 g10129(.a(new_n3058), .O(new_n10323));
  nor2 g10130(.a(new_n10320), .b(new_n2184), .O(new_n10324));
  inv1 g10131(.a(new_n10324), .O(new_n10325));
  nor2 g10132(.a(new_n10325), .b(new_n10323), .O(new_n10326));
  nor2 g10133(.a(new_n10326), .b(new_n10322), .O(new_n10327));
  nor2 g10134(.a(new_n10327), .b(new_n10319), .O(new_n10328));
  inv1 g10135(.a(new_n10327), .O(new_n10329));
  nor2 g10136(.a(new_n10329), .b(new_n10318), .O(new_n10330));
  nor2 g10137(.a(new_n10330), .b(new_n10328), .O(new_n10331));
  inv1 g10138(.a(new_n10331), .O(new_n10332));
  nor2 g10139(.a(new_n4425), .b(new_n1297), .O(new_n10333));
  nor2 g10140(.a(new_n4093), .b(new_n1493), .O(new_n10334));
  nor2 g10141(.a(new_n10334), .b(new_n9865), .O(new_n10335));
  inv1 g10142(.a(new_n9862), .O(new_n10336));
  nor2 g10143(.a(new_n4366), .b(new_n1493), .O(new_n10337));
  inv1 g10144(.a(new_n10337), .O(new_n10338));
  nor2 g10145(.a(new_n10338), .b(new_n10336), .O(new_n10339));
  nor2 g10146(.a(new_n10339), .b(new_n10335), .O(new_n10340));
  inv1 g10147(.a(new_n10340), .O(new_n10341));
  nor2 g10148(.a(new_n10341), .b(new_n10333), .O(new_n10342));
  inv1 g10149(.a(new_n10333), .O(new_n10343));
  nor2 g10150(.a(new_n10340), .b(new_n10343), .O(new_n10344));
  nor2 g10151(.a(new_n10344), .b(new_n10342), .O(new_n10345));
  nor2 g10152(.a(new_n3870), .b(new_n1647), .O(new_n10346));
  inv1 g10153(.a(new_n10346), .O(new_n10347));
  nor2 g10154(.a(new_n3533), .b(new_n1903), .O(new_n10348));
  nor2 g10155(.a(new_n10348), .b(new_n9925), .O(new_n10349));
  inv1 g10156(.a(new_n9923), .O(new_n10350));
  nor2 g10157(.a(new_n3722), .b(new_n1903), .O(new_n10351));
  inv1 g10158(.a(new_n10351), .O(new_n10352));
  nor2 g10159(.a(new_n10352), .b(new_n10350), .O(new_n10353));
  nor2 g10160(.a(new_n10353), .b(new_n10349), .O(new_n10354));
  nor2 g10161(.a(new_n10354), .b(new_n10347), .O(new_n10355));
  inv1 g10162(.a(new_n10354), .O(new_n10356));
  nor2 g10163(.a(new_n10356), .b(new_n10346), .O(new_n10357));
  nor2 g10164(.a(new_n10357), .b(new_n10355), .O(new_n10358));
  nor2 g10165(.a(new_n10358), .b(new_n10345), .O(new_n10359));
  inv1 g10166(.a(new_n10345), .O(new_n10360));
  inv1 g10167(.a(new_n10358), .O(new_n10361));
  nor2 g10168(.a(new_n10361), .b(new_n10360), .O(new_n10362));
  nor2 g10169(.a(new_n10362), .b(new_n10359), .O(new_n10363));
  nor2 g10170(.a(new_n10363), .b(new_n10332), .O(new_n10364));
  inv1 g10171(.a(new_n10363), .O(new_n10365));
  nor2 g10172(.a(new_n10365), .b(new_n10331), .O(new_n10366));
  nor2 g10173(.a(new_n10366), .b(new_n10364), .O(new_n10367));
  inv1 g10174(.a(new_n10367), .O(new_n10368));
  nor2 g10175(.a(new_n10368), .b(new_n10317), .O(new_n10369));
  nor2 g10176(.a(new_n10367), .b(new_n10316), .O(new_n10370));
  nor2 g10177(.a(new_n10370), .b(new_n10369), .O(new_n10371));
  inv1 g10178(.a(new_n10371), .O(new_n10372));
  nor2 g10179(.a(new_n10372), .b(new_n10272), .O(new_n10373));
  nor2 g10180(.a(new_n10371), .b(new_n10271), .O(new_n10374));
  nor2 g10181(.a(new_n10374), .b(new_n10373), .O(new_n10375));
  inv1 g10182(.a(new_n10375), .O(new_n10376));
  nor2 g10183(.a(new_n10376), .b(new_n10175), .O(new_n10377));
  nor2 g10184(.a(new_n10375), .b(new_n10174), .O(new_n10378));
  nor2 g10185(.a(new_n10378), .b(new_n10377), .O(new_n10379));
  inv1 g10186(.a(new_n10379), .O(new_n10380));
  nor2 g10187(.a(new_n10380), .b(new_n10092), .O(new_n10381));
  nor2 g10188(.a(new_n10379), .b(new_n10091), .O(new_n10382));
  nor2 g10189(.a(new_n10382), .b(new_n10381), .O(new_n10383));
  nor2 g10190(.a(new_n10035), .b(new_n9761), .O(new_n10384));
  inv1 g10191(.a(new_n10384), .O(new_n10385));
  nor2 g10192(.a(new_n10385), .b(new_n10383), .O(new_n10386));
  inv1 g10193(.a(new_n10383), .O(new_n10387));
  nor2 g10194(.a(new_n10384), .b(new_n10387), .O(new_n10388));
  nor2 g10195(.a(new_n10388), .b(new_n10386), .O(new_n10389));
  inv1 g10196(.a(new_n10389), .O(new_n10390));
  nor2 g10197(.a(new_n10044), .b(new_n10040), .O(new_n10391));
  nor2 g10198(.a(new_n10391), .b(new_n10390), .O(new_n10392));
  inv1 g10199(.a(new_n10391), .O(new_n10393));
  nor2 g10200(.a(new_n10393), .b(new_n10389), .O(new_n10394));
  nor2 g10201(.a(new_n10394), .b(new_n10392), .O(new_n10395));
  inv1 g10202(.a(new_n10395), .O(\asquared[60] ));
  nor2 g10203(.a(new_n10381), .b(new_n10090), .O(new_n10397));
  inv1 g10204(.a(new_n10397), .O(new_n10398));
  nor2 g10205(.a(new_n10377), .b(new_n10171), .O(new_n10399));
  inv1 g10206(.a(new_n10399), .O(new_n10400));
  nor2 g10207(.a(new_n10373), .b(new_n10270), .O(new_n10401));
  nor2 g10208(.a(new_n10167), .b(new_n10162), .O(new_n10402));
  nor2 g10209(.a(new_n10134), .b(new_n10128), .O(new_n10403));
  inv1 g10210(.a(new_n10403), .O(new_n10404));
  nor2 g10211(.a(new_n10120), .b(new_n10114), .O(new_n10405));
  inv1 g10212(.a(new_n10405), .O(new_n10406));
  nor2 g10213(.a(new_n10406), .b(new_n10404), .O(new_n10407));
  nor2 g10214(.a(new_n10405), .b(new_n10403), .O(new_n10408));
  nor2 g10215(.a(new_n10408), .b(new_n10407), .O(new_n10409));
  nor2 g10216(.a(new_n10209), .b(new_n10204), .O(new_n10410));
  inv1 g10217(.a(new_n10410), .O(new_n10411));
  nor2 g10218(.a(new_n10411), .b(new_n10409), .O(new_n10412));
  inv1 g10219(.a(new_n10409), .O(new_n10413));
  nor2 g10220(.a(new_n10410), .b(new_n10413), .O(new_n10414));
  nor2 g10221(.a(new_n10414), .b(new_n10412), .O(new_n10415));
  nor2 g10222(.a(new_n10105), .b(new_n10099), .O(new_n10416));
  inv1 g10223(.a(new_n10416), .O(new_n10417));
  nor2 g10224(.a(new_n10417), .b(new_n10415), .O(new_n10418));
  inv1 g10225(.a(new_n10415), .O(new_n10419));
  nor2 g10226(.a(new_n10416), .b(new_n10419), .O(new_n10420));
  nor2 g10227(.a(new_n10420), .b(new_n10418), .O(new_n10421));
  inv1 g10228(.a(new_n10421), .O(new_n10422));
  nor2 g10229(.a(new_n10369), .b(new_n10315), .O(new_n10423));
  nor2 g10230(.a(new_n10423), .b(new_n10422), .O(new_n10424));
  inv1 g10231(.a(new_n10423), .O(new_n10425));
  nor2 g10232(.a(new_n10425), .b(new_n10421), .O(new_n10426));
  nor2 g10233(.a(new_n10426), .b(new_n10424), .O(new_n10427));
  inv1 g10234(.a(new_n10427), .O(new_n10428));
  nor2 g10235(.a(new_n10428), .b(new_n10402), .O(new_n10429));
  inv1 g10236(.a(new_n10402), .O(new_n10430));
  nor2 g10237(.a(new_n10427), .b(new_n10430), .O(new_n10431));
  nor2 g10238(.a(new_n10431), .b(new_n10429), .O(new_n10432));
  inv1 g10239(.a(new_n10432), .O(new_n10433));
  nor2 g10240(.a(new_n10433), .b(new_n10401), .O(new_n10434));
  inv1 g10241(.a(new_n10401), .O(new_n10435));
  nor2 g10242(.a(new_n10432), .b(new_n10435), .O(new_n10436));
  nor2 g10243(.a(new_n10436), .b(new_n10434), .O(new_n10437));
  nor2 g10244(.a(new_n10437), .b(new_n10400), .O(new_n10438));
  inv1 g10245(.a(new_n10437), .O(new_n10439));
  nor2 g10246(.a(new_n10439), .b(new_n10399), .O(new_n10440));
  nor2 g10247(.a(new_n10440), .b(new_n10438), .O(new_n10441));
  inv1 g10248(.a(new_n10441), .O(new_n10442));
  nor2 g10249(.a(new_n10158), .b(new_n10154), .O(new_n10443));
  nor2 g10250(.a(new_n10150), .b(new_n10145), .O(new_n10444));
  inv1 g10251(.a(new_n10444), .O(new_n10445));
  nor2 g10252(.a(new_n3231), .b(new_n2184), .O(new_n10446));
  inv1 g10253(.a(new_n10446), .O(new_n10447));
  nor2 g10254(.a(new_n3057), .b(new_n2433), .O(new_n10448));
  nor2 g10255(.a(new_n4093), .b(new_n1647), .O(new_n10449));
  nor2 g10256(.a(new_n10449), .b(new_n10448), .O(new_n10450));
  inv1 g10257(.a(new_n10448), .O(new_n10451));
  inv1 g10258(.a(new_n10449), .O(new_n10452));
  nor2 g10259(.a(new_n10452), .b(new_n10451), .O(new_n10453));
  nor2 g10260(.a(new_n10453), .b(new_n10450), .O(new_n10454));
  nor2 g10261(.a(new_n10454), .b(new_n10447), .O(new_n10455));
  inv1 g10262(.a(new_n10454), .O(new_n10456));
  nor2 g10263(.a(new_n10456), .b(new_n10446), .O(new_n10457));
  nor2 g10264(.a(new_n10457), .b(new_n10455), .O(new_n10458));
  nor2 g10265(.a(new_n2826), .b(new_n2506), .O(new_n10459));
  nor2 g10266(.a(new_n10320), .b(new_n194), .O(new_n10460));
  nor2 g10267(.a(new_n10460), .b(new_n10459), .O(new_n10461));
  inv1 g10268(.a(new_n10459), .O(new_n10462));
  inv1 g10269(.a(new_n10460), .O(new_n10463));
  nor2 g10270(.a(new_n10463), .b(new_n10462), .O(new_n10464));
  nor2 g10271(.a(new_n10464), .b(new_n10461), .O(new_n10465));
  inv1 g10272(.a(new_n10465), .O(new_n10466));
  inv1 g10273(.a(new_n10137), .O(new_n10467));
  inv1 g10274(.a(\a[60] ), .O(new_n10468));
  nor2 g10275(.a(new_n10468), .b(new_n198), .O(new_n10469));
  inv1 g10276(.a(new_n10469), .O(new_n10470));
  nor2 g10277(.a(new_n10470), .b(new_n10467), .O(new_n10471));
  nor2 g10278(.a(new_n10469), .b(new_n10137), .O(new_n10472));
  nor2 g10279(.a(new_n10472), .b(new_n10471), .O(new_n10473));
  inv1 g10280(.a(new_n10473), .O(new_n10474));
  nor2 g10281(.a(new_n10474), .b(new_n10466), .O(new_n10475));
  nor2 g10282(.a(new_n10473), .b(new_n10465), .O(new_n10476));
  nor2 g10283(.a(new_n10476), .b(new_n10475), .O(new_n10477));
  inv1 g10284(.a(new_n10477), .O(new_n10478));
  nor2 g10285(.a(new_n10478), .b(new_n10458), .O(new_n10479));
  inv1 g10286(.a(new_n10458), .O(new_n10480));
  nor2 g10287(.a(new_n10477), .b(new_n10480), .O(new_n10481));
  nor2 g10288(.a(new_n10481), .b(new_n10479), .O(new_n10482));
  nor2 g10289(.a(new_n10482), .b(new_n10445), .O(new_n10483));
  inv1 g10290(.a(new_n10482), .O(new_n10484));
  nor2 g10291(.a(new_n10484), .b(new_n10444), .O(new_n10485));
  nor2 g10292(.a(new_n10485), .b(new_n10483), .O(new_n10486));
  nor2 g10293(.a(new_n8946), .b(new_n229), .O(new_n10487));
  inv1 g10294(.a(new_n10487), .O(new_n10488));
  nor2 g10295(.a(new_n8476), .b(new_n257), .O(new_n10489));
  nor2 g10296(.a(new_n4954), .b(new_n1199), .O(new_n10490));
  nor2 g10297(.a(new_n10490), .b(new_n10489), .O(new_n10491));
  inv1 g10298(.a(new_n10489), .O(new_n10492));
  inv1 g10299(.a(new_n10490), .O(new_n10493));
  nor2 g10300(.a(new_n10493), .b(new_n10492), .O(new_n10494));
  nor2 g10301(.a(new_n10494), .b(new_n10491), .O(new_n10495));
  nor2 g10302(.a(new_n10495), .b(new_n10488), .O(new_n10496));
  inv1 g10303(.a(new_n10495), .O(new_n10497));
  nor2 g10304(.a(new_n10497), .b(new_n10487), .O(new_n10498));
  nor2 g10305(.a(new_n10498), .b(new_n10496), .O(new_n10499));
  inv1 g10306(.a(new_n10499), .O(new_n10500));
  nor2 g10307(.a(new_n6893), .b(new_n569), .O(new_n10501));
  nor2 g10308(.a(new_n6570), .b(new_n613), .O(new_n10502));
  nor2 g10309(.a(new_n10502), .b(new_n10501), .O(new_n10503));
  inv1 g10310(.a(new_n10227), .O(new_n10504));
  nor2 g10311(.a(new_n6893), .b(new_n613), .O(new_n10505));
  inv1 g10312(.a(new_n10505), .O(new_n10506));
  nor2 g10313(.a(new_n10506), .b(new_n10504), .O(new_n10507));
  nor2 g10314(.a(new_n10507), .b(new_n10503), .O(new_n10508));
  nor2 g10315(.a(new_n10508), .b(new_n9110), .O(new_n10509));
  inv1 g10316(.a(new_n10508), .O(new_n10510));
  nor2 g10317(.a(new_n10510), .b(new_n9109), .O(new_n10511));
  nor2 g10318(.a(new_n10511), .b(new_n10509), .O(new_n10512));
  nor2 g10319(.a(new_n8170), .b(new_n295), .O(new_n10513));
  inv1 g10320(.a(new_n10513), .O(new_n10514));
  nor2 g10321(.a(new_n8026), .b(new_n322), .O(new_n10515));
  nor2 g10322(.a(new_n5178), .b(new_n1086), .O(new_n10516));
  nor2 g10323(.a(new_n10516), .b(new_n10515), .O(new_n10517));
  inv1 g10324(.a(new_n10515), .O(new_n10518));
  inv1 g10325(.a(new_n10516), .O(new_n10519));
  nor2 g10326(.a(new_n10519), .b(new_n10518), .O(new_n10520));
  nor2 g10327(.a(new_n10520), .b(new_n10517), .O(new_n10521));
  nor2 g10328(.a(new_n10521), .b(new_n10514), .O(new_n10522));
  inv1 g10329(.a(new_n10521), .O(new_n10523));
  nor2 g10330(.a(new_n10523), .b(new_n10513), .O(new_n10524));
  nor2 g10331(.a(new_n10524), .b(new_n10522), .O(new_n10525));
  nor2 g10332(.a(new_n10525), .b(new_n10512), .O(new_n10526));
  inv1 g10333(.a(new_n10512), .O(new_n10527));
  inv1 g10334(.a(new_n10525), .O(new_n10528));
  nor2 g10335(.a(new_n10528), .b(new_n10527), .O(new_n10529));
  nor2 g10336(.a(new_n10529), .b(new_n10526), .O(new_n10530));
  nor2 g10337(.a(new_n10530), .b(new_n10500), .O(new_n10531));
  inv1 g10338(.a(new_n10530), .O(new_n10532));
  nor2 g10339(.a(new_n10532), .b(new_n10499), .O(new_n10533));
  nor2 g10340(.a(new_n10533), .b(new_n10531), .O(new_n10534));
  nor2 g10341(.a(new_n10534), .b(new_n10486), .O(new_n10535));
  inv1 g10342(.a(new_n10486), .O(new_n10536));
  inv1 g10343(.a(new_n10534), .O(new_n10537));
  nor2 g10344(.a(new_n10537), .b(new_n10536), .O(new_n10538));
  nor2 g10345(.a(new_n10538), .b(new_n10535), .O(new_n10539));
  inv1 g10346(.a(new_n10539), .O(new_n10540));
  nor2 g10347(.a(new_n10540), .b(new_n10443), .O(new_n10541));
  inv1 g10348(.a(new_n10443), .O(new_n10542));
  nor2 g10349(.a(new_n10539), .b(new_n10542), .O(new_n10543));
  nor2 g10350(.a(new_n10543), .b(new_n10541), .O(new_n10544));
  inv1 g10351(.a(new_n10544), .O(new_n10545));
  nor2 g10352(.a(new_n10074), .b(new_n10069), .O(new_n10546));
  nor2 g10353(.a(new_n10065), .b(new_n10059), .O(new_n10547));
  inv1 g10354(.a(new_n10547), .O(new_n10548));
  nor2 g10355(.a(new_n3870), .b(new_n1736), .O(new_n10549));
  inv1 g10356(.a(new_n10549), .O(new_n10550));
  nor2 g10357(.a(new_n3533), .b(new_n2121), .O(new_n10551));
  nor2 g10358(.a(new_n10551), .b(new_n10351), .O(new_n10552));
  inv1 g10359(.a(new_n10348), .O(new_n10553));
  nor2 g10360(.a(new_n3722), .b(new_n2121), .O(new_n10554));
  inv1 g10361(.a(new_n10554), .O(new_n10555));
  nor2 g10362(.a(new_n10555), .b(new_n10553), .O(new_n10556));
  nor2 g10363(.a(new_n10556), .b(new_n10552), .O(new_n10557));
  nor2 g10364(.a(new_n10557), .b(new_n10550), .O(new_n10558));
  inv1 g10365(.a(new_n10557), .O(new_n10559));
  nor2 g10366(.a(new_n10559), .b(new_n10549), .O(new_n10560));
  nor2 g10367(.a(new_n10560), .b(new_n10558), .O(new_n10561));
  inv1 g10368(.a(new_n10561), .O(new_n10562));
  nor2 g10369(.a(new_n9873), .b(new_n196), .O(new_n10563));
  nor2 g10370(.a(new_n9156), .b(new_n214), .O(new_n10564));
  nor2 g10371(.a(new_n10564), .b(new_n10193), .O(new_n10565));
  inv1 g10372(.a(new_n10191), .O(new_n10566));
  nor2 g10373(.a(new_n9658), .b(new_n214), .O(new_n10567));
  inv1 g10374(.a(new_n10567), .O(new_n10568));
  nor2 g10375(.a(new_n10568), .b(new_n10566), .O(new_n10569));
  nor2 g10376(.a(new_n10569), .b(new_n10565), .O(new_n10570));
  inv1 g10377(.a(new_n10570), .O(new_n10571));
  nor2 g10378(.a(new_n10571), .b(new_n10563), .O(new_n10572));
  inv1 g10379(.a(new_n10563), .O(new_n10573));
  nor2 g10380(.a(new_n10570), .b(new_n10573), .O(new_n10574));
  nor2 g10381(.a(new_n10574), .b(new_n10572), .O(new_n10575));
  nor2 g10382(.a(new_n4682), .b(new_n1297), .O(new_n10576));
  inv1 g10383(.a(new_n10576), .O(new_n10577));
  nor2 g10384(.a(new_n4425), .b(new_n1425), .O(new_n10578));
  nor2 g10385(.a(new_n10578), .b(new_n10337), .O(new_n10579));
  nor2 g10386(.a(new_n4425), .b(new_n1493), .O(new_n10580));
  inv1 g10387(.a(new_n10580), .O(new_n10581));
  nor2 g10388(.a(new_n10581), .b(new_n9866), .O(new_n10582));
  nor2 g10389(.a(new_n10582), .b(new_n10579), .O(new_n10583));
  nor2 g10390(.a(new_n10583), .b(new_n10577), .O(new_n10584));
  inv1 g10391(.a(new_n10583), .O(new_n10585));
  nor2 g10392(.a(new_n10585), .b(new_n10576), .O(new_n10586));
  nor2 g10393(.a(new_n10586), .b(new_n10584), .O(new_n10587));
  nor2 g10394(.a(new_n10587), .b(new_n10575), .O(new_n10588));
  inv1 g10395(.a(new_n10575), .O(new_n10589));
  inv1 g10396(.a(new_n10587), .O(new_n10590));
  nor2 g10397(.a(new_n10590), .b(new_n10589), .O(new_n10591));
  nor2 g10398(.a(new_n10591), .b(new_n10588), .O(new_n10592));
  nor2 g10399(.a(new_n10592), .b(new_n10562), .O(new_n10593));
  inv1 g10400(.a(new_n10592), .O(new_n10594));
  nor2 g10401(.a(new_n10594), .b(new_n10561), .O(new_n10595));
  nor2 g10402(.a(new_n10595), .b(new_n10593), .O(new_n10596));
  nor2 g10403(.a(new_n10596), .b(new_n10548), .O(new_n10597));
  inv1 g10404(.a(new_n10596), .O(new_n10598));
  nor2 g10405(.a(new_n10598), .b(new_n10547), .O(new_n10599));
  nor2 g10406(.a(new_n10599), .b(new_n10597), .O(new_n10600));
  nor2 g10407(.a(new_n7294), .b(new_n438), .O(new_n10601));
  inv1 g10408(.a(new_n10601), .O(new_n10602));
  nor2 g10409(.a(new_n6958), .b(new_n502), .O(new_n10603));
  nor2 g10410(.a(new_n10603), .b(new_n7237), .O(new_n10604));
  nor2 g10411(.a(new_n10295), .b(new_n9072), .O(new_n10605));
  nor2 g10412(.a(new_n10605), .b(new_n10604), .O(new_n10606));
  nor2 g10413(.a(new_n10606), .b(new_n10602), .O(new_n10607));
  inv1 g10414(.a(new_n10606), .O(new_n10608));
  nor2 g10415(.a(new_n10608), .b(new_n10601), .O(new_n10609));
  nor2 g10416(.a(new_n10609), .b(new_n10607), .O(new_n10610));
  nor2 g10417(.a(new_n7537), .b(new_n363), .O(new_n10611));
  nor2 g10418(.a(new_n5796), .b(new_n847), .O(new_n10612));
  nor2 g10419(.a(new_n10612), .b(new_n10611), .O(new_n10613));
  inv1 g10420(.a(new_n8197), .O(new_n10614));
  nor2 g10421(.a(new_n7537), .b(new_n847), .O(new_n10615));
  inv1 g10422(.a(new_n10615), .O(new_n10616));
  nor2 g10423(.a(new_n10616), .b(new_n10614), .O(new_n10617));
  nor2 g10424(.a(new_n10617), .b(new_n10613), .O(new_n10618));
  nor2 g10425(.a(new_n10618), .b(new_n10218), .O(new_n10619));
  inv1 g10426(.a(new_n10618), .O(new_n10620));
  nor2 g10427(.a(new_n10620), .b(new_n10217), .O(new_n10621));
  nor2 g10428(.a(new_n10621), .b(new_n10619), .O(new_n10622));
  nor2 g10429(.a(new_n10234), .b(new_n10228), .O(new_n10623));
  inv1 g10430(.a(new_n10623), .O(new_n10624));
  nor2 g10431(.a(new_n10624), .b(new_n10622), .O(new_n10625));
  inv1 g10432(.a(new_n10622), .O(new_n10626));
  nor2 g10433(.a(new_n10623), .b(new_n10626), .O(new_n10627));
  nor2 g10434(.a(new_n10627), .b(new_n10625), .O(new_n10628));
  inv1 g10435(.a(new_n10628), .O(new_n10629));
  nor2 g10436(.a(new_n10629), .b(new_n10610), .O(new_n10630));
  inv1 g10437(.a(new_n10610), .O(new_n10631));
  nor2 g10438(.a(new_n10628), .b(new_n10631), .O(new_n10632));
  nor2 g10439(.a(new_n10632), .b(new_n10630), .O(new_n10633));
  nor2 g10440(.a(new_n10633), .b(new_n10600), .O(new_n10634));
  inv1 g10441(.a(new_n10600), .O(new_n10635));
  inv1 g10442(.a(new_n10633), .O(new_n10636));
  nor2 g10443(.a(new_n10636), .b(new_n10635), .O(new_n10637));
  nor2 g10444(.a(new_n10637), .b(new_n10634), .O(new_n10638));
  inv1 g10445(.a(new_n10638), .O(new_n10639));
  nor2 g10446(.a(new_n10639), .b(new_n10546), .O(new_n10640));
  inv1 g10447(.a(new_n10546), .O(new_n10641));
  nor2 g10448(.a(new_n10638), .b(new_n10641), .O(new_n10642));
  nor2 g10449(.a(new_n10642), .b(new_n10640), .O(new_n10643));
  inv1 g10450(.a(new_n10643), .O(new_n10644));
  nor2 g10451(.a(new_n10644), .b(new_n10545), .O(new_n10645));
  nor2 g10452(.a(new_n10643), .b(new_n10544), .O(new_n10646));
  nor2 g10453(.a(new_n10646), .b(new_n10645), .O(new_n10647));
  inv1 g10454(.a(new_n10647), .O(new_n10648));
  nor2 g10455(.a(new_n10084), .b(new_n10079), .O(new_n10649));
  nor2 g10456(.a(new_n10223), .b(new_n10215), .O(new_n10650));
  nor2 g10457(.a(new_n10284), .b(new_n10278), .O(new_n10651));
  nor2 g10458(.a(new_n10651), .b(new_n10650), .O(new_n10652));
  inv1 g10459(.a(new_n10650), .O(new_n10653));
  inv1 g10460(.a(new_n10651), .O(new_n10654));
  nor2 g10461(.a(new_n10654), .b(new_n10653), .O(new_n10655));
  nor2 g10462(.a(new_n10655), .b(new_n10652), .O(new_n10656));
  nor2 g10463(.a(new_n10247), .b(new_n10240), .O(new_n10657));
  nor2 g10464(.a(new_n10657), .b(new_n10656), .O(new_n10658));
  inv1 g10465(.a(new_n10656), .O(new_n10659));
  inv1 g10466(.a(new_n10657), .O(new_n10660));
  nor2 g10467(.a(new_n10660), .b(new_n10659), .O(new_n10661));
  nor2 g10468(.a(new_n10661), .b(new_n10658), .O(new_n10662));
  nor2 g10469(.a(new_n10366), .b(new_n10359), .O(new_n10663));
  inv1 g10470(.a(new_n10663), .O(new_n10664));
  nor2 g10471(.a(new_n10664), .b(new_n10662), .O(new_n10665));
  inv1 g10472(.a(new_n10662), .O(new_n10666));
  nor2 g10473(.a(new_n10663), .b(new_n10666), .O(new_n10667));
  nor2 g10474(.a(new_n10667), .b(new_n10665), .O(new_n10668));
  nor2 g10475(.a(new_n10256), .b(new_n10249), .O(new_n10669));
  inv1 g10476(.a(new_n10669), .O(new_n10670));
  nor2 g10477(.a(new_n10670), .b(new_n10668), .O(new_n10671));
  inv1 g10478(.a(new_n10668), .O(new_n10672));
  nor2 g10479(.a(new_n10669), .b(new_n10672), .O(new_n10673));
  nor2 g10480(.a(new_n10673), .b(new_n10671), .O(new_n10674));
  inv1 g10481(.a(new_n10674), .O(new_n10675));
  nor2 g10482(.a(new_n10264), .b(new_n10261), .O(new_n10676));
  nor2 g10483(.a(new_n10309), .b(new_n10302), .O(new_n10677));
  nor2 g10484(.a(new_n10188), .b(new_n10181), .O(new_n10678));
  nor2 g10485(.a(new_n10342), .b(new_n10335), .O(new_n10679));
  nor2 g10486(.a(new_n10679), .b(new_n10678), .O(new_n10680));
  inv1 g10487(.a(new_n10678), .O(new_n10681));
  inv1 g10488(.a(new_n10679), .O(new_n10682));
  nor2 g10489(.a(new_n10682), .b(new_n10681), .O(new_n10683));
  nor2 g10490(.a(new_n10683), .b(new_n10680), .O(new_n10684));
  nor2 g10491(.a(new_n10357), .b(new_n10349), .O(new_n10685));
  nor2 g10492(.a(new_n10685), .b(new_n10684), .O(new_n10686));
  inv1 g10493(.a(new_n10684), .O(new_n10687));
  inv1 g10494(.a(new_n10685), .O(new_n10688));
  nor2 g10495(.a(new_n10688), .b(new_n10687), .O(new_n10689));
  nor2 g10496(.a(new_n10689), .b(new_n10686), .O(new_n10690));
  inv1 g10497(.a(new_n10690), .O(new_n10691));
  nor2 g10498(.a(new_n10330), .b(new_n10322), .O(new_n10692));
  nor2 g10499(.a(new_n10198), .b(new_n10192), .O(new_n10693));
  nor2 g10500(.a(new_n10693), .b(new_n10692), .O(new_n10694));
  inv1 g10501(.a(new_n10692), .O(new_n10695));
  inv1 g10502(.a(new_n10693), .O(new_n10696));
  nor2 g10503(.a(new_n10696), .b(new_n10695), .O(new_n10697));
  nor2 g10504(.a(new_n10697), .b(new_n10694), .O(new_n10698));
  nor2 g10505(.a(new_n10300), .b(new_n10292), .O(new_n10699));
  nor2 g10506(.a(new_n10699), .b(new_n10698), .O(new_n10700));
  inv1 g10507(.a(new_n10698), .O(new_n10701));
  inv1 g10508(.a(new_n10699), .O(new_n10702));
  nor2 g10509(.a(new_n10702), .b(new_n10701), .O(new_n10703));
  nor2 g10510(.a(new_n10703), .b(new_n10700), .O(new_n10704));
  inv1 g10511(.a(new_n10704), .O(new_n10705));
  nor2 g10512(.a(new_n10705), .b(new_n10691), .O(new_n10706));
  nor2 g10513(.a(new_n10704), .b(new_n10690), .O(new_n10707));
  nor2 g10514(.a(new_n10707), .b(new_n10706), .O(new_n10708));
  inv1 g10515(.a(new_n10708), .O(new_n10709));
  nor2 g10516(.a(new_n10709), .b(new_n10677), .O(new_n10710));
  inv1 g10517(.a(new_n10677), .O(new_n10711));
  nor2 g10518(.a(new_n10708), .b(new_n10711), .O(new_n10712));
  nor2 g10519(.a(new_n10712), .b(new_n10710), .O(new_n10713));
  inv1 g10520(.a(new_n10713), .O(new_n10714));
  nor2 g10521(.a(new_n10714), .b(new_n10676), .O(new_n10715));
  inv1 g10522(.a(new_n10676), .O(new_n10716));
  nor2 g10523(.a(new_n10713), .b(new_n10716), .O(new_n10717));
  nor2 g10524(.a(new_n10717), .b(new_n10715), .O(new_n10718));
  inv1 g10525(.a(new_n10718), .O(new_n10719));
  nor2 g10526(.a(new_n10719), .b(new_n10675), .O(new_n10720));
  nor2 g10527(.a(new_n10718), .b(new_n10674), .O(new_n10721));
  nor2 g10528(.a(new_n10721), .b(new_n10720), .O(new_n10722));
  inv1 g10529(.a(new_n10722), .O(new_n10723));
  nor2 g10530(.a(new_n10723), .b(new_n10649), .O(new_n10724));
  inv1 g10531(.a(new_n10649), .O(new_n10725));
  nor2 g10532(.a(new_n10722), .b(new_n10725), .O(new_n10726));
  nor2 g10533(.a(new_n10726), .b(new_n10724), .O(new_n10727));
  inv1 g10534(.a(new_n10727), .O(new_n10728));
  nor2 g10535(.a(new_n10728), .b(new_n10648), .O(new_n10729));
  nor2 g10536(.a(new_n10727), .b(new_n10647), .O(new_n10730));
  nor2 g10537(.a(new_n10730), .b(new_n10729), .O(new_n10731));
  inv1 g10538(.a(new_n10731), .O(new_n10732));
  nor2 g10539(.a(new_n10732), .b(new_n10442), .O(new_n10733));
  nor2 g10540(.a(new_n10731), .b(new_n10441), .O(new_n10734));
  nor2 g10541(.a(new_n10734), .b(new_n10733), .O(new_n10735));
  nor2 g10542(.a(new_n10735), .b(new_n10398), .O(new_n10736));
  inv1 g10543(.a(new_n10735), .O(new_n10737));
  nor2 g10544(.a(new_n10737), .b(new_n10397), .O(new_n10738));
  nor2 g10545(.a(new_n10738), .b(new_n10736), .O(new_n10739));
  inv1 g10546(.a(new_n10739), .O(new_n10740));
  nor2 g10547(.a(new_n10392), .b(new_n10386), .O(new_n10741));
  nor2 g10548(.a(new_n10741), .b(new_n10740), .O(new_n10742));
  inv1 g10549(.a(new_n10741), .O(new_n10743));
  nor2 g10550(.a(new_n10743), .b(new_n10739), .O(new_n10744));
  nor2 g10551(.a(new_n10744), .b(new_n10742), .O(new_n10745));
  inv1 g10552(.a(new_n10745), .O(\asquared[61] ));
  nor2 g10553(.a(new_n10733), .b(new_n10440), .O(new_n10747));
  nor2 g10554(.a(new_n10434), .b(new_n10429), .O(new_n10748));
  inv1 g10555(.a(new_n10748), .O(new_n10749));
  nor2 g10556(.a(new_n10541), .b(new_n10538), .O(new_n10750));
  inv1 g10557(.a(new_n10750), .O(new_n10751));
  nor2 g10558(.a(new_n10524), .b(new_n10517), .O(new_n10752));
  nor2 g10559(.a(new_n10621), .b(new_n10613), .O(new_n10753));
  nor2 g10560(.a(new_n10753), .b(new_n10752), .O(new_n10754));
  inv1 g10561(.a(new_n10752), .O(new_n10755));
  inv1 g10562(.a(new_n10753), .O(new_n10756));
  nor2 g10563(.a(new_n10756), .b(new_n10755), .O(new_n10757));
  nor2 g10564(.a(new_n10757), .b(new_n10754), .O(new_n10758));
  nor2 g10565(.a(new_n10475), .b(new_n10471), .O(new_n10759));
  inv1 g10566(.a(new_n10759), .O(new_n10760));
  nor2 g10567(.a(new_n10760), .b(new_n10758), .O(new_n10761));
  inv1 g10568(.a(new_n10758), .O(new_n10762));
  nor2 g10569(.a(new_n10759), .b(new_n10762), .O(new_n10763));
  nor2 g10570(.a(new_n10763), .b(new_n10761), .O(new_n10764));
  nor2 g10571(.a(new_n10533), .b(new_n10526), .O(new_n10765));
  inv1 g10572(.a(new_n10765), .O(new_n10766));
  nor2 g10573(.a(new_n10766), .b(new_n10764), .O(new_n10767));
  inv1 g10574(.a(new_n10764), .O(new_n10768));
  nor2 g10575(.a(new_n10765), .b(new_n10768), .O(new_n10769));
  nor2 g10576(.a(new_n10769), .b(new_n10767), .O(new_n10770));
  nor2 g10577(.a(new_n10485), .b(new_n10479), .O(new_n10771));
  inv1 g10578(.a(new_n10771), .O(new_n10772));
  nor2 g10579(.a(new_n10772), .b(new_n10770), .O(new_n10773));
  inv1 g10580(.a(new_n10770), .O(new_n10774));
  nor2 g10581(.a(new_n10771), .b(new_n10774), .O(new_n10775));
  nor2 g10582(.a(new_n10775), .b(new_n10773), .O(new_n10776));
  nor2 g10583(.a(new_n10457), .b(new_n10450), .O(new_n10777));
  nor2 g10584(.a(new_n10560), .b(new_n10552), .O(new_n10778));
  nor2 g10585(.a(new_n10778), .b(new_n10777), .O(new_n10779));
  inv1 g10586(.a(new_n10777), .O(new_n10780));
  inv1 g10587(.a(new_n10778), .O(new_n10781));
  nor2 g10588(.a(new_n10781), .b(new_n10780), .O(new_n10782));
  nor2 g10589(.a(new_n10782), .b(new_n10779), .O(new_n10783));
  nor2 g10590(.a(new_n10586), .b(new_n10579), .O(new_n10784));
  nor2 g10591(.a(new_n10784), .b(new_n10783), .O(new_n10785));
  inv1 g10592(.a(new_n10783), .O(new_n10786));
  inv1 g10593(.a(new_n10784), .O(new_n10787));
  nor2 g10594(.a(new_n10787), .b(new_n10786), .O(new_n10788));
  nor2 g10595(.a(new_n10788), .b(new_n10785), .O(new_n10789));
  nor2 g10596(.a(new_n10498), .b(new_n10491), .O(new_n10790));
  nor2 g10597(.a(new_n10572), .b(new_n10565), .O(new_n10791));
  nor2 g10598(.a(new_n10791), .b(new_n10790), .O(new_n10792));
  inv1 g10599(.a(new_n10790), .O(new_n10793));
  inv1 g10600(.a(new_n10791), .O(new_n10794));
  nor2 g10601(.a(new_n10794), .b(new_n10793), .O(new_n10795));
  nor2 g10602(.a(new_n10795), .b(new_n10792), .O(new_n10796));
  nor2 g10603(.a(new_n10609), .b(new_n10604), .O(new_n10797));
  nor2 g10604(.a(new_n10797), .b(new_n10796), .O(new_n10798));
  inv1 g10605(.a(new_n10796), .O(new_n10799));
  inv1 g10606(.a(new_n10797), .O(new_n10800));
  nor2 g10607(.a(new_n10800), .b(new_n10799), .O(new_n10801));
  nor2 g10608(.a(new_n10801), .b(new_n10798), .O(new_n10802));
  nor2 g10609(.a(new_n10802), .b(new_n10789), .O(new_n10803));
  inv1 g10610(.a(new_n10789), .O(new_n10804));
  inv1 g10611(.a(new_n10802), .O(new_n10805));
  nor2 g10612(.a(new_n10805), .b(new_n10804), .O(new_n10806));
  nor2 g10613(.a(new_n10806), .b(new_n10803), .O(new_n10807));
  inv1 g10614(.a(new_n10807), .O(new_n10808));
  nor2 g10615(.a(new_n10595), .b(new_n10588), .O(new_n10809));
  nor2 g10616(.a(new_n10809), .b(new_n10808), .O(new_n10810));
  inv1 g10617(.a(new_n10809), .O(new_n10811));
  nor2 g10618(.a(new_n10811), .b(new_n10807), .O(new_n10812));
  nor2 g10619(.a(new_n10812), .b(new_n10810), .O(new_n10813));
  nor2 g10620(.a(new_n10813), .b(new_n10776), .O(new_n10814));
  inv1 g10621(.a(new_n10776), .O(new_n10815));
  inv1 g10622(.a(new_n10813), .O(new_n10816));
  nor2 g10623(.a(new_n10816), .b(new_n10815), .O(new_n10817));
  nor2 g10624(.a(new_n10817), .b(new_n10814), .O(new_n10818));
  inv1 g10625(.a(new_n10818), .O(new_n10819));
  nor2 g10626(.a(new_n10819), .b(new_n10751), .O(new_n10820));
  nor2 g10627(.a(new_n10818), .b(new_n10750), .O(new_n10821));
  nor2 g10628(.a(new_n10821), .b(new_n10820), .O(new_n10822));
  inv1 g10629(.a(new_n10822), .O(new_n10823));
  nor2 g10630(.a(new_n10823), .b(new_n10749), .O(new_n10824));
  nor2 g10631(.a(new_n10822), .b(new_n10748), .O(new_n10825));
  nor2 g10632(.a(new_n10825), .b(new_n10824), .O(new_n10826));
  inv1 g10633(.a(new_n10826), .O(new_n10827));
  nor2 g10634(.a(new_n10720), .b(new_n10715), .O(new_n10828));
  nor2 g10635(.a(new_n10424), .b(new_n10420), .O(new_n10829));
  nor2 g10636(.a(new_n10414), .b(new_n10408), .O(new_n10830));
  inv1 g10637(.a(new_n10830), .O(new_n10831));
  nor2 g10638(.a(new_n2826), .b(new_n2660), .O(new_n10832));
  nor2 g10639(.a(new_n3057), .b(new_n2506), .O(new_n10833));
  nor2 g10640(.a(new_n10833), .b(new_n10832), .O(new_n10834));
  nor2 g10641(.a(new_n3057), .b(new_n2660), .O(new_n10835));
  inv1 g10642(.a(new_n10835), .O(new_n10836));
  nor2 g10643(.a(new_n10836), .b(new_n10462), .O(new_n10837));
  nor2 g10644(.a(new_n10837), .b(new_n10834), .O(new_n10838));
  nor2 g10645(.a(new_n10838), .b(new_n10506), .O(new_n10839));
  inv1 g10646(.a(new_n10838), .O(new_n10840));
  nor2 g10647(.a(new_n10840), .b(new_n10505), .O(new_n10841));
  nor2 g10648(.a(new_n10841), .b(new_n10839), .O(new_n10842));
  nor2 g10649(.a(new_n7294), .b(new_n502), .O(new_n10843));
  inv1 g10650(.a(new_n10843), .O(new_n10844));
  nor2 g10651(.a(new_n6958), .b(new_n569), .O(new_n10845));
  nor2 g10652(.a(new_n10845), .b(new_n10229), .O(new_n10846));
  nor2 g10653(.a(new_n6958), .b(new_n699), .O(new_n10847));
  inv1 g10654(.a(new_n10847), .O(new_n10848));
  nor2 g10655(.a(new_n10848), .b(new_n10504), .O(new_n10849));
  nor2 g10656(.a(new_n10849), .b(new_n10846), .O(new_n10850));
  nor2 g10657(.a(new_n10850), .b(new_n10844), .O(new_n10851));
  inv1 g10658(.a(new_n10850), .O(new_n10852));
  nor2 g10659(.a(new_n10852), .b(new_n10843), .O(new_n10853));
  nor2 g10660(.a(new_n10853), .b(new_n10851), .O(new_n10854));
  nor2 g10661(.a(new_n5971), .b(new_n847), .O(new_n10855));
  inv1 g10662(.a(new_n10855), .O(new_n10856));
  nor2 g10663(.a(new_n6274), .b(new_n800), .O(new_n10857));
  nor2 g10664(.a(new_n7537), .b(new_n438), .O(new_n10858));
  nor2 g10665(.a(new_n10858), .b(new_n10857), .O(new_n10859));
  inv1 g10666(.a(new_n9107), .O(new_n10860));
  nor2 g10667(.a(new_n7537), .b(new_n800), .O(new_n10861));
  inv1 g10668(.a(new_n10861), .O(new_n10862));
  nor2 g10669(.a(new_n10862), .b(new_n10860), .O(new_n10863));
  nor2 g10670(.a(new_n10863), .b(new_n10859), .O(new_n10864));
  nor2 g10671(.a(new_n10864), .b(new_n10856), .O(new_n10865));
  inv1 g10672(.a(new_n10864), .O(new_n10866));
  nor2 g10673(.a(new_n10866), .b(new_n10855), .O(new_n10867));
  nor2 g10674(.a(new_n10867), .b(new_n10865), .O(new_n10868));
  nor2 g10675(.a(new_n10868), .b(new_n10854), .O(new_n10869));
  inv1 g10676(.a(new_n10854), .O(new_n10870));
  inv1 g10677(.a(new_n10868), .O(new_n10871));
  nor2 g10678(.a(new_n10871), .b(new_n10870), .O(new_n10872));
  nor2 g10679(.a(new_n10872), .b(new_n10869), .O(new_n10873));
  inv1 g10680(.a(new_n10873), .O(new_n10874));
  nor2 g10681(.a(new_n10874), .b(new_n10842), .O(new_n10875));
  inv1 g10682(.a(new_n10842), .O(new_n10876));
  nor2 g10683(.a(new_n10873), .b(new_n10876), .O(new_n10877));
  nor2 g10684(.a(new_n10877), .b(new_n10875), .O(new_n10878));
  nor2 g10685(.a(new_n10878), .b(new_n10831), .O(new_n10879));
  inv1 g10686(.a(new_n10878), .O(new_n10880));
  nor2 g10687(.a(new_n10880), .b(new_n10830), .O(new_n10881));
  nor2 g10688(.a(new_n10881), .b(new_n10879), .O(new_n10882));
  nor2 g10689(.a(new_n4093), .b(new_n1736), .O(new_n10883));
  nor2 g10690(.a(new_n3870), .b(new_n1903), .O(new_n10884));
  nor2 g10691(.a(new_n10884), .b(new_n10883), .O(new_n10885));
  nor2 g10692(.a(new_n4093), .b(new_n1903), .O(new_n10886));
  inv1 g10693(.a(new_n10886), .O(new_n10887));
  nor2 g10694(.a(new_n10887), .b(new_n10550), .O(new_n10888));
  nor2 g10695(.a(new_n10888), .b(new_n10885), .O(new_n10889));
  nor2 g10696(.a(new_n10889), .b(new_n10581), .O(new_n10890));
  inv1 g10697(.a(new_n10889), .O(new_n10891));
  nor2 g10698(.a(new_n10891), .b(new_n10580), .O(new_n10892));
  nor2 g10699(.a(new_n10892), .b(new_n10890), .O(new_n10893));
  inv1 g10700(.a(new_n10893), .O(new_n10894));
  inv1 g10701(.a(\a[61] ), .O(new_n10895));
  nor2 g10702(.a(new_n10895), .b(new_n198), .O(new_n10896));
  nor2 g10703(.a(new_n10320), .b(new_n196), .O(new_n10897));
  nor2 g10704(.a(new_n9156), .b(new_n229), .O(new_n10898));
  nor2 g10705(.a(new_n10898), .b(new_n10897), .O(new_n10899));
  nor2 g10706(.a(new_n10320), .b(new_n229), .O(new_n10900));
  inv1 g10707(.a(new_n10900), .O(new_n10901));
  nor2 g10708(.a(new_n10901), .b(new_n9161), .O(new_n10902));
  nor2 g10709(.a(new_n10902), .b(new_n10899), .O(new_n10903));
  inv1 g10710(.a(new_n10903), .O(new_n10904));
  nor2 g10711(.a(new_n10904), .b(new_n10896), .O(new_n10905));
  inv1 g10712(.a(new_n10896), .O(new_n10906));
  nor2 g10713(.a(new_n10903), .b(new_n10906), .O(new_n10907));
  nor2 g10714(.a(new_n10907), .b(new_n10905), .O(new_n10908));
  nor2 g10715(.a(new_n8946), .b(new_n257), .O(new_n10909));
  inv1 g10716(.a(new_n10909), .O(new_n10910));
  nor2 g10717(.a(new_n4954), .b(new_n1297), .O(new_n10911));
  nor2 g10718(.a(new_n4682), .b(new_n1425), .O(new_n10912));
  nor2 g10719(.a(new_n10912), .b(new_n10911), .O(new_n10913));
  nor2 g10720(.a(new_n4954), .b(new_n1425), .O(new_n10914));
  inv1 g10721(.a(new_n10914), .O(new_n10915));
  nor2 g10722(.a(new_n10915), .b(new_n10577), .O(new_n10916));
  nor2 g10723(.a(new_n10916), .b(new_n10913), .O(new_n10917));
  nor2 g10724(.a(new_n10917), .b(new_n10910), .O(new_n10918));
  inv1 g10725(.a(new_n10917), .O(new_n10919));
  nor2 g10726(.a(new_n10919), .b(new_n10909), .O(new_n10920));
  nor2 g10727(.a(new_n10920), .b(new_n10918), .O(new_n10921));
  nor2 g10728(.a(new_n10921), .b(new_n10908), .O(new_n10922));
  inv1 g10729(.a(new_n10908), .O(new_n10923));
  inv1 g10730(.a(new_n10921), .O(new_n10924));
  nor2 g10731(.a(new_n10924), .b(new_n10923), .O(new_n10925));
  nor2 g10732(.a(new_n10925), .b(new_n10922), .O(new_n10926));
  nor2 g10733(.a(new_n10926), .b(new_n10894), .O(new_n10927));
  inv1 g10734(.a(new_n10926), .O(new_n10928));
  nor2 g10735(.a(new_n10928), .b(new_n10893), .O(new_n10929));
  nor2 g10736(.a(new_n10929), .b(new_n10927), .O(new_n10930));
  nor2 g10737(.a(new_n10930), .b(new_n10882), .O(new_n10931));
  inv1 g10738(.a(new_n10882), .O(new_n10932));
  inv1 g10739(.a(new_n10930), .O(new_n10933));
  nor2 g10740(.a(new_n10933), .b(new_n10932), .O(new_n10934));
  nor2 g10741(.a(new_n10934), .b(new_n10931), .O(new_n10935));
  inv1 g10742(.a(new_n10935), .O(new_n10936));
  nor2 g10743(.a(new_n10936), .b(new_n10829), .O(new_n10937));
  inv1 g10744(.a(new_n10829), .O(new_n10938));
  nor2 g10745(.a(new_n10935), .b(new_n10938), .O(new_n10939));
  nor2 g10746(.a(new_n10939), .b(new_n10937), .O(new_n10940));
  inv1 g10747(.a(new_n10940), .O(new_n10941));
  nor2 g10748(.a(new_n10941), .b(new_n10828), .O(new_n10942));
  inv1 g10749(.a(new_n10828), .O(new_n10943));
  nor2 g10750(.a(new_n10940), .b(new_n10943), .O(new_n10944));
  nor2 g10751(.a(new_n10944), .b(new_n10942), .O(new_n10945));
  inv1 g10752(.a(new_n10945), .O(new_n10946));
  nor2 g10753(.a(new_n10946), .b(new_n10827), .O(new_n10947));
  nor2 g10754(.a(new_n10945), .b(new_n10826), .O(new_n10948));
  nor2 g10755(.a(new_n10948), .b(new_n10947), .O(new_n10949));
  inv1 g10756(.a(new_n10949), .O(new_n10950));
  nor2 g10757(.a(new_n10729), .b(new_n10724), .O(new_n10951));
  nor2 g10758(.a(new_n10645), .b(new_n10640), .O(new_n10952));
  nor2 g10759(.a(new_n10637), .b(new_n10599), .O(new_n10953));
  nor2 g10760(.a(new_n10630), .b(new_n10625), .O(new_n10954));
  nor2 g10761(.a(new_n10689), .b(new_n10683), .O(new_n10955));
  nor2 g10762(.a(new_n10468), .b(new_n194), .O(new_n10956));
  inv1 g10763(.a(new_n10956), .O(new_n10957));
  nor2 g10764(.a(new_n10464), .b(new_n2826), .O(new_n10958));
  nor2 g10765(.a(new_n10958), .b(new_n10957), .O(new_n10959));
  inv1 g10766(.a(new_n10958), .O(new_n10960));
  nor2 g10767(.a(new_n10960), .b(new_n10956), .O(new_n10961));
  nor2 g10768(.a(new_n10961), .b(new_n10959), .O(new_n10962));
  nor2 g10769(.a(new_n10511), .b(new_n10503), .O(new_n10963));
  inv1 g10770(.a(new_n10963), .O(new_n10964));
  nor2 g10771(.a(new_n10964), .b(new_n10962), .O(new_n10965));
  inv1 g10772(.a(new_n10962), .O(new_n10966));
  nor2 g10773(.a(new_n10963), .b(new_n10966), .O(new_n10967));
  nor2 g10774(.a(new_n10967), .b(new_n10965), .O(new_n10968));
  inv1 g10775(.a(new_n10968), .O(new_n10969));
  nor2 g10776(.a(new_n10969), .b(new_n10955), .O(new_n10970));
  inv1 g10777(.a(new_n10955), .O(new_n10971));
  nor2 g10778(.a(new_n10968), .b(new_n10971), .O(new_n10972));
  nor2 g10779(.a(new_n10972), .b(new_n10970), .O(new_n10973));
  inv1 g10780(.a(new_n10973), .O(new_n10974));
  nor2 g10781(.a(new_n10974), .b(new_n10954), .O(new_n10975));
  inv1 g10782(.a(new_n10954), .O(new_n10976));
  nor2 g10783(.a(new_n10973), .b(new_n10976), .O(new_n10977));
  nor2 g10784(.a(new_n10977), .b(new_n10975), .O(new_n10978));
  inv1 g10785(.a(new_n10978), .O(new_n10979));
  nor2 g10786(.a(new_n10703), .b(new_n10697), .O(new_n10980));
  nor2 g10787(.a(new_n10661), .b(new_n10655), .O(new_n10981));
  nor2 g10788(.a(new_n4366), .b(new_n1647), .O(new_n10982));
  inv1 g10789(.a(new_n10982), .O(new_n10983));
  nor2 g10790(.a(new_n9873), .b(new_n203), .O(new_n10984));
  nor2 g10791(.a(new_n10984), .b(new_n10567), .O(new_n10985));
  nor2 g10792(.a(new_n9873), .b(new_n214), .O(new_n10986));
  inv1 g10793(.a(new_n10986), .O(new_n10987));
  nor2 g10794(.a(new_n10987), .b(new_n10194), .O(new_n10988));
  nor2 g10795(.a(new_n10988), .b(new_n10985), .O(new_n10989));
  nor2 g10796(.a(new_n10989), .b(new_n10983), .O(new_n10990));
  inv1 g10797(.a(new_n10989), .O(new_n10991));
  nor2 g10798(.a(new_n10991), .b(new_n10982), .O(new_n10992));
  nor2 g10799(.a(new_n10992), .b(new_n10990), .O(new_n10993));
  nor2 g10800(.a(new_n10993), .b(new_n10981), .O(new_n10994));
  inv1 g10801(.a(new_n10981), .O(new_n10995));
  inv1 g10802(.a(new_n10993), .O(new_n10996));
  nor2 g10803(.a(new_n10996), .b(new_n10995), .O(new_n10997));
  nor2 g10804(.a(new_n10997), .b(new_n10994), .O(new_n10998));
  inv1 g10805(.a(new_n10998), .O(new_n10999));
  nor2 g10806(.a(new_n10999), .b(new_n10980), .O(new_n11000));
  inv1 g10807(.a(new_n10980), .O(new_n11001));
  nor2 g10808(.a(new_n10998), .b(new_n11001), .O(new_n11002));
  nor2 g10809(.a(new_n11002), .b(new_n11000), .O(new_n11003));
  inv1 g10810(.a(new_n11003), .O(new_n11004));
  nor2 g10811(.a(new_n11004), .b(new_n10979), .O(new_n11005));
  nor2 g10812(.a(new_n11003), .b(new_n10978), .O(new_n11006));
  nor2 g10813(.a(new_n11006), .b(new_n11005), .O(new_n11007));
  inv1 g10814(.a(new_n11007), .O(new_n11008));
  nor2 g10815(.a(new_n11008), .b(new_n10953), .O(new_n11009));
  inv1 g10816(.a(new_n10953), .O(new_n11010));
  nor2 g10817(.a(new_n11007), .b(new_n11010), .O(new_n11011));
  nor2 g10818(.a(new_n11011), .b(new_n11009), .O(new_n11012));
  inv1 g10819(.a(new_n11012), .O(new_n11013));
  nor2 g10820(.a(new_n10673), .b(new_n10667), .O(new_n11014));
  nor2 g10821(.a(new_n10710), .b(new_n10706), .O(new_n11015));
  nor2 g10822(.a(new_n3533), .b(new_n2184), .O(new_n11016));
  nor2 g10823(.a(new_n3231), .b(new_n2433), .O(new_n11017));
  nor2 g10824(.a(new_n11017), .b(new_n11016), .O(new_n11018));
  nor2 g10825(.a(new_n3533), .b(new_n2433), .O(new_n11019));
  inv1 g10826(.a(new_n11019), .O(new_n11020));
  nor2 g10827(.a(new_n11020), .b(new_n10447), .O(new_n11021));
  nor2 g10828(.a(new_n11021), .b(new_n11018), .O(new_n11022));
  nor2 g10829(.a(new_n11022), .b(new_n10555), .O(new_n11023));
  inv1 g10830(.a(new_n11022), .O(new_n11024));
  nor2 g10831(.a(new_n11024), .b(new_n10554), .O(new_n11025));
  nor2 g10832(.a(new_n11025), .b(new_n11023), .O(new_n11026));
  inv1 g10833(.a(new_n11026), .O(new_n11027));
  nor2 g10834(.a(new_n5178), .b(new_n1199), .O(new_n11028));
  nor2 g10835(.a(new_n8476), .b(new_n295), .O(new_n11029));
  nor2 g10836(.a(new_n8170), .b(new_n322), .O(new_n11030));
  nor2 g10837(.a(new_n11030), .b(new_n11029), .O(new_n11031));
  nor2 g10838(.a(new_n8476), .b(new_n322), .O(new_n11032));
  inv1 g10839(.a(new_n11032), .O(new_n11033));
  nor2 g10840(.a(new_n11033), .b(new_n10514), .O(new_n11034));
  nor2 g10841(.a(new_n11034), .b(new_n11031), .O(new_n11035));
  inv1 g10842(.a(new_n11035), .O(new_n11036));
  nor2 g10843(.a(new_n11036), .b(new_n11028), .O(new_n11037));
  inv1 g10844(.a(new_n11028), .O(new_n11038));
  nor2 g10845(.a(new_n11035), .b(new_n11038), .O(new_n11039));
  nor2 g10846(.a(new_n11039), .b(new_n11037), .O(new_n11040));
  nor2 g10847(.a(new_n5393), .b(new_n1086), .O(new_n11041));
  inv1 g10848(.a(new_n11041), .O(new_n11042));
  nor2 g10849(.a(new_n8026), .b(new_n363), .O(new_n11043));
  nor2 g10850(.a(new_n5796), .b(new_n941), .O(new_n11044));
  nor2 g10851(.a(new_n11044), .b(new_n11043), .O(new_n11045));
  nor2 g10852(.a(new_n8026), .b(new_n941), .O(new_n11046));
  inv1 g10853(.a(new_n11046), .O(new_n11047));
  nor2 g10854(.a(new_n11047), .b(new_n10614), .O(new_n11048));
  nor2 g10855(.a(new_n11048), .b(new_n11045), .O(new_n11049));
  nor2 g10856(.a(new_n11049), .b(new_n11042), .O(new_n11050));
  inv1 g10857(.a(new_n11049), .O(new_n11051));
  nor2 g10858(.a(new_n11051), .b(new_n11041), .O(new_n11052));
  nor2 g10859(.a(new_n11052), .b(new_n11050), .O(new_n11053));
  nor2 g10860(.a(new_n11053), .b(new_n11040), .O(new_n11054));
  inv1 g10861(.a(new_n11040), .O(new_n11055));
  inv1 g10862(.a(new_n11053), .O(new_n11056));
  nor2 g10863(.a(new_n11056), .b(new_n11055), .O(new_n11057));
  nor2 g10864(.a(new_n11057), .b(new_n11054), .O(new_n11058));
  nor2 g10865(.a(new_n11058), .b(new_n11027), .O(new_n11059));
  inv1 g10866(.a(new_n11058), .O(new_n11060));
  nor2 g10867(.a(new_n11060), .b(new_n11026), .O(new_n11061));
  nor2 g10868(.a(new_n11061), .b(new_n11059), .O(new_n11062));
  inv1 g10869(.a(new_n11062), .O(new_n11063));
  nor2 g10870(.a(new_n11063), .b(new_n11015), .O(new_n11064));
  inv1 g10871(.a(new_n11015), .O(new_n11065));
  nor2 g10872(.a(new_n11062), .b(new_n11065), .O(new_n11066));
  nor2 g10873(.a(new_n11066), .b(new_n11064), .O(new_n11067));
  inv1 g10874(.a(new_n11067), .O(new_n11068));
  nor2 g10875(.a(new_n11068), .b(new_n11014), .O(new_n11069));
  inv1 g10876(.a(new_n11014), .O(new_n11070));
  nor2 g10877(.a(new_n11067), .b(new_n11070), .O(new_n11071));
  nor2 g10878(.a(new_n11071), .b(new_n11069), .O(new_n11072));
  inv1 g10879(.a(new_n11072), .O(new_n11073));
  nor2 g10880(.a(new_n11073), .b(new_n11013), .O(new_n11074));
  nor2 g10881(.a(new_n11072), .b(new_n11012), .O(new_n11075));
  nor2 g10882(.a(new_n11075), .b(new_n11074), .O(new_n11076));
  inv1 g10883(.a(new_n11076), .O(new_n11077));
  nor2 g10884(.a(new_n11077), .b(new_n10952), .O(new_n11078));
  inv1 g10885(.a(new_n10952), .O(new_n11079));
  nor2 g10886(.a(new_n11076), .b(new_n11079), .O(new_n11080));
  nor2 g10887(.a(new_n11080), .b(new_n11078), .O(new_n11081));
  inv1 g10888(.a(new_n11081), .O(new_n11082));
  nor2 g10889(.a(new_n11082), .b(new_n10951), .O(new_n11083));
  inv1 g10890(.a(new_n10951), .O(new_n11084));
  nor2 g10891(.a(new_n11081), .b(new_n11084), .O(new_n11085));
  nor2 g10892(.a(new_n11085), .b(new_n11083), .O(new_n11086));
  inv1 g10893(.a(new_n11086), .O(new_n11087));
  nor2 g10894(.a(new_n11087), .b(new_n10950), .O(new_n11088));
  nor2 g10895(.a(new_n11086), .b(new_n10949), .O(new_n11089));
  nor2 g10896(.a(new_n11089), .b(new_n11088), .O(new_n11090));
  inv1 g10897(.a(new_n11090), .O(new_n11091));
  nor2 g10898(.a(new_n11091), .b(new_n10747), .O(new_n11092));
  inv1 g10899(.a(new_n10747), .O(new_n11093));
  nor2 g10900(.a(new_n11090), .b(new_n11093), .O(new_n11094));
  nor2 g10901(.a(new_n11094), .b(new_n11092), .O(new_n11095));
  inv1 g10902(.a(new_n11095), .O(new_n11096));
  nor2 g10903(.a(new_n10742), .b(new_n10736), .O(new_n11097));
  nor2 g10904(.a(new_n11097), .b(new_n11096), .O(new_n11098));
  inv1 g10905(.a(new_n11097), .O(new_n11099));
  nor2 g10906(.a(new_n11099), .b(new_n11095), .O(new_n11100));
  nor2 g10907(.a(new_n11100), .b(new_n11098), .O(new_n11101));
  inv1 g10908(.a(new_n11101), .O(\asquared[62] ));
  nor2 g10909(.a(new_n11088), .b(new_n11083), .O(new_n11103));
  nor2 g10910(.a(new_n11078), .b(new_n11074), .O(new_n11104));
  nor2 g10911(.a(new_n11052), .b(new_n11045), .O(new_n11105));
  nor2 g10912(.a(new_n10867), .b(new_n10859), .O(new_n11106));
  nor2 g10913(.a(new_n11106), .b(new_n11105), .O(new_n11107));
  inv1 g10914(.a(new_n11105), .O(new_n11108));
  inv1 g10915(.a(new_n11106), .O(new_n11109));
  nor2 g10916(.a(new_n11109), .b(new_n11108), .O(new_n11110));
  nor2 g10917(.a(new_n11110), .b(new_n11107), .O(new_n11111));
  inv1 g10918(.a(new_n11111), .O(new_n11112));
  nor2 g10919(.a(new_n10320), .b(new_n203), .O(new_n11113));
  inv1 g10920(.a(new_n11113), .O(new_n11114));
  nor2 g10921(.a(new_n9658), .b(new_n229), .O(new_n11115));
  nor2 g10922(.a(new_n11115), .b(new_n10986), .O(new_n11116));
  nor2 g10923(.a(new_n9873), .b(new_n229), .O(new_n11117));
  inv1 g10924(.a(new_n11117), .O(new_n11118));
  nor2 g10925(.a(new_n11118), .b(new_n10568), .O(new_n11119));
  nor2 g10926(.a(new_n11119), .b(new_n11116), .O(new_n11120));
  nor2 g10927(.a(new_n11120), .b(new_n11114), .O(new_n11121));
  inv1 g10928(.a(new_n11120), .O(new_n11122));
  nor2 g10929(.a(new_n11122), .b(new_n11113), .O(new_n11123));
  nor2 g10930(.a(new_n11123), .b(new_n11121), .O(new_n11124));
  nor2 g10931(.a(new_n11124), .b(new_n11112), .O(new_n11125));
  inv1 g10932(.a(new_n11124), .O(new_n11126));
  nor2 g10933(.a(new_n11126), .b(new_n11111), .O(new_n11127));
  nor2 g10934(.a(new_n11127), .b(new_n11125), .O(new_n11128));
  nor2 g10935(.a(new_n11061), .b(new_n11054), .O(new_n11129));
  inv1 g10936(.a(new_n11129), .O(new_n11130));
  nor2 g10937(.a(new_n11130), .b(new_n11128), .O(new_n11131));
  inv1 g10938(.a(new_n11128), .O(new_n11132));
  nor2 g10939(.a(new_n11129), .b(new_n11132), .O(new_n11133));
  nor2 g10940(.a(new_n11133), .b(new_n11131), .O(new_n11134));
  nor2 g10941(.a(new_n11000), .b(new_n10994), .O(new_n11135));
  inv1 g10942(.a(new_n11135), .O(new_n11136));
  nor2 g10943(.a(new_n11136), .b(new_n11134), .O(new_n11137));
  inv1 g10944(.a(new_n11134), .O(new_n11138));
  nor2 g10945(.a(new_n11135), .b(new_n11138), .O(new_n11139));
  nor2 g10946(.a(new_n11139), .b(new_n11137), .O(new_n11140));
  inv1 g10947(.a(new_n11140), .O(new_n11141));
  nor2 g10948(.a(new_n10763), .b(new_n10757), .O(new_n11142));
  inv1 g10949(.a(new_n11142), .O(new_n11143));
  inv1 g10950(.a(new_n10464), .O(new_n11144));
  nor2 g10951(.a(new_n11144), .b(\a[60] ), .O(new_n11145));
  nor2 g10952(.a(new_n11145), .b(new_n10965), .O(new_n11146));
  inv1 g10953(.a(new_n11146), .O(new_n11147));
  nor2 g10954(.a(new_n11147), .b(new_n11143), .O(new_n11148));
  nor2 g10955(.a(new_n11146), .b(new_n11142), .O(new_n11149));
  nor2 g10956(.a(new_n11149), .b(new_n11148), .O(new_n11150));
  nor2 g10957(.a(new_n10788), .b(new_n10782), .O(new_n11151));
  inv1 g10958(.a(new_n11151), .O(new_n11152));
  nor2 g10959(.a(new_n11152), .b(new_n11150), .O(new_n11153));
  inv1 g10960(.a(new_n11150), .O(new_n11154));
  nor2 g10961(.a(new_n11151), .b(new_n11154), .O(new_n11155));
  nor2 g10962(.a(new_n11155), .b(new_n11153), .O(new_n11156));
  inv1 g10963(.a(new_n11156), .O(new_n11157));
  nor2 g10964(.a(new_n10934), .b(new_n10881), .O(new_n11158));
  nor2 g10965(.a(new_n11158), .b(new_n11157), .O(new_n11159));
  inv1 g10966(.a(new_n11158), .O(new_n11160));
  nor2 g10967(.a(new_n11160), .b(new_n11156), .O(new_n11161));
  nor2 g10968(.a(new_n11161), .b(new_n11159), .O(new_n11162));
  inv1 g10969(.a(new_n11162), .O(new_n11163));
  nor2 g10970(.a(new_n11163), .b(new_n11141), .O(new_n11164));
  nor2 g10971(.a(new_n11162), .b(new_n11140), .O(new_n11165));
  nor2 g10972(.a(new_n11165), .b(new_n11164), .O(new_n11166));
  inv1 g10973(.a(new_n11166), .O(new_n11167));
  nor2 g10974(.a(new_n11167), .b(new_n11104), .O(new_n11168));
  inv1 g10975(.a(new_n11104), .O(new_n11169));
  nor2 g10976(.a(new_n11166), .b(new_n11169), .O(new_n11170));
  nor2 g10977(.a(new_n11170), .b(new_n11168), .O(new_n11171));
  nor2 g10978(.a(new_n11009), .b(new_n11005), .O(new_n11172));
  nor2 g10979(.a(new_n8170), .b(new_n363), .O(new_n11173));
  inv1 g10980(.a(new_n11173), .O(new_n11174));
  nor2 g10981(.a(new_n8026), .b(new_n438), .O(new_n11175));
  nor2 g10982(.a(new_n5971), .b(new_n941), .O(new_n11176));
  nor2 g10983(.a(new_n11176), .b(new_n11175), .O(new_n11177));
  nor2 g10984(.a(new_n11047), .b(new_n8886), .O(new_n11178));
  nor2 g10985(.a(new_n11178), .b(new_n11177), .O(new_n11179));
  nor2 g10986(.a(new_n11179), .b(new_n11174), .O(new_n11180));
  inv1 g10987(.a(new_n11179), .O(new_n11181));
  nor2 g10988(.a(new_n11181), .b(new_n11173), .O(new_n11182));
  nor2 g10989(.a(new_n11182), .b(new_n11180), .O(new_n11183));
  inv1 g10990(.a(new_n11183), .O(new_n11184));
  nor2 g10991(.a(new_n10957), .b(new_n2826), .O(new_n11185));
  inv1 g10992(.a(\a[62] ), .O(new_n11186));
  nor2 g10993(.a(new_n11186), .b(new_n198), .O(new_n11187));
  nor2 g10994(.a(new_n10468), .b(new_n196), .O(new_n11188));
  nor2 g10995(.a(new_n11188), .b(new_n11187), .O(new_n11189));
  nor2 g10996(.a(new_n11186), .b(new_n196), .O(new_n11190));
  inv1 g10997(.a(new_n11190), .O(new_n11191));
  nor2 g10998(.a(new_n11191), .b(new_n10470), .O(new_n11192));
  nor2 g10999(.a(new_n11192), .b(new_n11189), .O(new_n11193));
  inv1 g11000(.a(new_n11193), .O(new_n11194));
  nor2 g11001(.a(new_n11194), .b(new_n11185), .O(new_n11195));
  inv1 g11002(.a(new_n11185), .O(new_n11196));
  nor2 g11003(.a(new_n11193), .b(new_n11196), .O(new_n11197));
  nor2 g11004(.a(new_n11197), .b(new_n11195), .O(new_n11198));
  nor2 g11005(.a(new_n3870), .b(new_n2121), .O(new_n11199));
  nor2 g11006(.a(new_n11199), .b(new_n10886), .O(new_n11200));
  inv1 g11007(.a(new_n10884), .O(new_n11201));
  nor2 g11008(.a(new_n4093), .b(new_n2121), .O(new_n11202));
  inv1 g11009(.a(new_n11202), .O(new_n11203));
  nor2 g11010(.a(new_n11203), .b(new_n11201), .O(new_n11204));
  nor2 g11011(.a(new_n11204), .b(new_n11200), .O(new_n11205));
  nor2 g11012(.a(new_n11205), .b(new_n10915), .O(new_n11206));
  inv1 g11013(.a(new_n11205), .O(new_n11207));
  nor2 g11014(.a(new_n11207), .b(new_n10914), .O(new_n11208));
  nor2 g11015(.a(new_n11208), .b(new_n11206), .O(new_n11209));
  nor2 g11016(.a(new_n11209), .b(new_n11198), .O(new_n11210));
  inv1 g11017(.a(new_n11198), .O(new_n11211));
  inv1 g11018(.a(new_n11209), .O(new_n11212));
  nor2 g11019(.a(new_n11212), .b(new_n11211), .O(new_n11213));
  nor2 g11020(.a(new_n11213), .b(new_n11210), .O(new_n11214));
  nor2 g11021(.a(new_n11214), .b(new_n11184), .O(new_n11215));
  inv1 g11022(.a(new_n11214), .O(new_n11216));
  nor2 g11023(.a(new_n11216), .b(new_n11183), .O(new_n11217));
  nor2 g11024(.a(new_n11217), .b(new_n11215), .O(new_n11218));
  inv1 g11025(.a(new_n11218), .O(new_n11219));
  nor2 g11026(.a(new_n5178), .b(new_n1297), .O(new_n11220));
  inv1 g11027(.a(new_n11220), .O(new_n11221));
  nor2 g11028(.a(new_n9156), .b(new_n257), .O(new_n11222));
  nor2 g11029(.a(new_n8946), .b(new_n295), .O(new_n11223));
  nor2 g11030(.a(new_n11223), .b(new_n11222), .O(new_n11224));
  nor2 g11031(.a(new_n9156), .b(new_n295), .O(new_n11225));
  inv1 g11032(.a(new_n11225), .O(new_n11226));
  nor2 g11033(.a(new_n11226), .b(new_n10910), .O(new_n11227));
  nor2 g11034(.a(new_n11227), .b(new_n11224), .O(new_n11228));
  nor2 g11035(.a(new_n11228), .b(new_n11221), .O(new_n11229));
  inv1 g11036(.a(new_n11228), .O(new_n11230));
  nor2 g11037(.a(new_n11230), .b(new_n11220), .O(new_n11231));
  nor2 g11038(.a(new_n11231), .b(new_n11229), .O(new_n11232));
  inv1 g11039(.a(new_n11232), .O(new_n11233));
  nor2 g11040(.a(new_n7537), .b(new_n502), .O(new_n11234));
  nor2 g11041(.a(new_n11234), .b(new_n9988), .O(new_n11235));
  inv1 g11042(.a(new_n9985), .O(new_n11236));
  nor2 g11043(.a(new_n10862), .b(new_n11236), .O(new_n11237));
  nor2 g11044(.a(new_n11237), .b(new_n11235), .O(new_n11238));
  inv1 g11045(.a(new_n11238), .O(new_n11239));
  nor2 g11046(.a(new_n11239), .b(new_n7853), .O(new_n11240));
  nor2 g11047(.a(new_n11238), .b(new_n7854), .O(new_n11241));
  nor2 g11048(.a(new_n11241), .b(new_n11240), .O(new_n11242));
  nor2 g11049(.a(new_n7294), .b(new_n569), .O(new_n11243));
  inv1 g11050(.a(new_n11243), .O(new_n11244));
  nor2 g11051(.a(new_n6958), .b(new_n613), .O(new_n11245));
  nor2 g11052(.a(new_n6893), .b(new_n699), .O(new_n11246));
  nor2 g11053(.a(new_n11246), .b(new_n11245), .O(new_n11247));
  nor2 g11054(.a(new_n10848), .b(new_n10506), .O(new_n11248));
  nor2 g11055(.a(new_n11248), .b(new_n11247), .O(new_n11249));
  nor2 g11056(.a(new_n11249), .b(new_n11244), .O(new_n11250));
  inv1 g11057(.a(new_n11249), .O(new_n11251));
  nor2 g11058(.a(new_n11251), .b(new_n11243), .O(new_n11252));
  nor2 g11059(.a(new_n11252), .b(new_n11250), .O(new_n11253));
  nor2 g11060(.a(new_n11253), .b(new_n11242), .O(new_n11254));
  inv1 g11061(.a(new_n11242), .O(new_n11255));
  inv1 g11062(.a(new_n11253), .O(new_n11256));
  nor2 g11063(.a(new_n11256), .b(new_n11255), .O(new_n11257));
  nor2 g11064(.a(new_n11257), .b(new_n11254), .O(new_n11258));
  nor2 g11065(.a(new_n11258), .b(new_n11233), .O(new_n11259));
  inv1 g11066(.a(new_n11258), .O(new_n11260));
  nor2 g11067(.a(new_n11260), .b(new_n11232), .O(new_n11261));
  nor2 g11068(.a(new_n11261), .b(new_n11259), .O(new_n11262));
  inv1 g11069(.a(new_n11262), .O(new_n11263));
  nor2 g11070(.a(new_n11263), .b(new_n11219), .O(new_n11264));
  nor2 g11071(.a(new_n11262), .b(new_n11218), .O(new_n11265));
  nor2 g11072(.a(new_n11265), .b(new_n11264), .O(new_n11266));
  inv1 g11073(.a(new_n11266), .O(new_n11267));
  nor2 g11074(.a(new_n4682), .b(new_n1493), .O(new_n11268));
  inv1 g11075(.a(new_n11268), .O(new_n11269));
  nor2 g11076(.a(new_n4425), .b(new_n1647), .O(new_n11270));
  nor2 g11077(.a(new_n4366), .b(new_n1736), .O(new_n11271));
  nor2 g11078(.a(new_n11271), .b(new_n11270), .O(new_n11272));
  nor2 g11079(.a(new_n4425), .b(new_n1736), .O(new_n11273));
  inv1 g11080(.a(new_n11273), .O(new_n11274));
  nor2 g11081(.a(new_n11274), .b(new_n10983), .O(new_n11275));
  nor2 g11082(.a(new_n11275), .b(new_n11272), .O(new_n11276));
  nor2 g11083(.a(new_n11276), .b(new_n11269), .O(new_n11277));
  inv1 g11084(.a(new_n11276), .O(new_n11278));
  nor2 g11085(.a(new_n11278), .b(new_n11268), .O(new_n11279));
  nor2 g11086(.a(new_n11279), .b(new_n11277), .O(new_n11280));
  inv1 g11087(.a(new_n11280), .O(new_n11281));
  nor2 g11088(.a(new_n5393), .b(new_n1199), .O(new_n11282));
  nor2 g11089(.a(new_n5796), .b(new_n1086), .O(new_n11283));
  nor2 g11090(.a(new_n11283), .b(new_n11032), .O(new_n11284));
  inv1 g11091(.a(new_n7828), .O(new_n11285));
  nor2 g11092(.a(new_n8476), .b(new_n1086), .O(new_n11286));
  inv1 g11093(.a(new_n11286), .O(new_n11287));
  nor2 g11094(.a(new_n11287), .b(new_n11285), .O(new_n11288));
  nor2 g11095(.a(new_n11288), .b(new_n11284), .O(new_n11289));
  inv1 g11096(.a(new_n11289), .O(new_n11290));
  nor2 g11097(.a(new_n11290), .b(new_n11282), .O(new_n11291));
  inv1 g11098(.a(new_n11282), .O(new_n11292));
  nor2 g11099(.a(new_n11289), .b(new_n11292), .O(new_n11293));
  nor2 g11100(.a(new_n11293), .b(new_n11291), .O(new_n11294));
  nor2 g11101(.a(new_n3722), .b(new_n2184), .O(new_n11295));
  inv1 g11102(.a(new_n11295), .O(new_n11296));
  nor2 g11103(.a(new_n3231), .b(new_n2506), .O(new_n11297));
  nor2 g11104(.a(new_n11297), .b(new_n11019), .O(new_n11298));
  inv1 g11105(.a(new_n11017), .O(new_n11299));
  nor2 g11106(.a(new_n3533), .b(new_n2506), .O(new_n11300));
  inv1 g11107(.a(new_n11300), .O(new_n11301));
  nor2 g11108(.a(new_n11301), .b(new_n11299), .O(new_n11302));
  nor2 g11109(.a(new_n11302), .b(new_n11298), .O(new_n11303));
  nor2 g11110(.a(new_n11303), .b(new_n11296), .O(new_n11304));
  inv1 g11111(.a(new_n11303), .O(new_n11305));
  nor2 g11112(.a(new_n11305), .b(new_n11295), .O(new_n11306));
  nor2 g11113(.a(new_n11306), .b(new_n11304), .O(new_n11307));
  nor2 g11114(.a(new_n11307), .b(new_n11294), .O(new_n11308));
  inv1 g11115(.a(new_n11294), .O(new_n11309));
  inv1 g11116(.a(new_n11307), .O(new_n11310));
  nor2 g11117(.a(new_n11310), .b(new_n11309), .O(new_n11311));
  nor2 g11118(.a(new_n11311), .b(new_n11308), .O(new_n11312));
  nor2 g11119(.a(new_n11312), .b(new_n11281), .O(new_n11313));
  inv1 g11120(.a(new_n11312), .O(new_n11314));
  nor2 g11121(.a(new_n11314), .b(new_n11280), .O(new_n11315));
  nor2 g11122(.a(new_n11315), .b(new_n11313), .O(new_n11316));
  inv1 g11123(.a(new_n11316), .O(new_n11317));
  nor2 g11124(.a(new_n11317), .b(new_n11267), .O(new_n11318));
  nor2 g11125(.a(new_n11316), .b(new_n11266), .O(new_n11319));
  nor2 g11126(.a(new_n11319), .b(new_n11318), .O(new_n11320));
  inv1 g11127(.a(new_n11320), .O(new_n11321));
  nor2 g11128(.a(new_n11321), .b(new_n11172), .O(new_n11322));
  inv1 g11129(.a(new_n11172), .O(new_n11323));
  nor2 g11130(.a(new_n11320), .b(new_n11323), .O(new_n11324));
  nor2 g11131(.a(new_n11324), .b(new_n11322), .O(new_n11325));
  inv1 g11132(.a(new_n11325), .O(new_n11326));
  nor2 g11133(.a(new_n10820), .b(new_n10814), .O(new_n11327));
  inv1 g11134(.a(new_n11327), .O(new_n11328));
  nor2 g11135(.a(new_n11328), .b(new_n11326), .O(new_n11329));
  nor2 g11136(.a(new_n11327), .b(new_n11325), .O(new_n11330));
  nor2 g11137(.a(new_n11330), .b(new_n11329), .O(new_n11331));
  nor2 g11138(.a(new_n11331), .b(new_n11171), .O(new_n11332));
  inv1 g11139(.a(new_n11171), .O(new_n11333));
  inv1 g11140(.a(new_n11331), .O(new_n11334));
  nor2 g11141(.a(new_n11334), .b(new_n11333), .O(new_n11335));
  nor2 g11142(.a(new_n11335), .b(new_n11332), .O(new_n11336));
  inv1 g11143(.a(new_n11336), .O(new_n11337));
  nor2 g11144(.a(new_n10947), .b(new_n10825), .O(new_n11338));
  nor2 g11145(.a(new_n11069), .b(new_n11064), .O(new_n11339));
  inv1 g11146(.a(new_n11339), .O(new_n11340));
  nor2 g11147(.a(new_n10801), .b(new_n10795), .O(new_n11341));
  inv1 g11148(.a(new_n11341), .O(new_n11342));
  nor2 g11149(.a(new_n10929), .b(new_n10922), .O(new_n11343));
  inv1 g11150(.a(new_n11343), .O(new_n11344));
  nor2 g11151(.a(new_n11344), .b(new_n11342), .O(new_n11345));
  nor2 g11152(.a(new_n11343), .b(new_n11341), .O(new_n11346));
  nor2 g11153(.a(new_n11346), .b(new_n11345), .O(new_n11347));
  nor2 g11154(.a(new_n10875), .b(new_n10869), .O(new_n11348));
  inv1 g11155(.a(new_n11348), .O(new_n11349));
  nor2 g11156(.a(new_n11349), .b(new_n11347), .O(new_n11350));
  inv1 g11157(.a(new_n11347), .O(new_n11351));
  nor2 g11158(.a(new_n11348), .b(new_n11351), .O(new_n11352));
  nor2 g11159(.a(new_n11352), .b(new_n11350), .O(new_n11353));
  inv1 g11160(.a(new_n11353), .O(new_n11354));
  nor2 g11161(.a(new_n10920), .b(new_n10913), .O(new_n11355));
  nor2 g11162(.a(new_n10905), .b(new_n10899), .O(new_n11356));
  nor2 g11163(.a(new_n11356), .b(new_n11355), .O(new_n11357));
  inv1 g11164(.a(new_n11355), .O(new_n11358));
  inv1 g11165(.a(new_n11356), .O(new_n11359));
  nor2 g11166(.a(new_n11359), .b(new_n11358), .O(new_n11360));
  nor2 g11167(.a(new_n11360), .b(new_n11357), .O(new_n11361));
  nor2 g11168(.a(new_n11037), .b(new_n11031), .O(new_n11362));
  nor2 g11169(.a(new_n11362), .b(new_n11361), .O(new_n11363));
  inv1 g11170(.a(new_n11361), .O(new_n11364));
  inv1 g11171(.a(new_n11362), .O(new_n11365));
  nor2 g11172(.a(new_n11365), .b(new_n11364), .O(new_n11366));
  nor2 g11173(.a(new_n11366), .b(new_n11363), .O(new_n11367));
  inv1 g11174(.a(new_n11367), .O(new_n11368));
  nor2 g11175(.a(new_n11025), .b(new_n11018), .O(new_n11369));
  nor2 g11176(.a(new_n10992), .b(new_n10985), .O(new_n11370));
  nor2 g11177(.a(new_n11370), .b(new_n11369), .O(new_n11371));
  inv1 g11178(.a(new_n11369), .O(new_n11372));
  inv1 g11179(.a(new_n11370), .O(new_n11373));
  nor2 g11180(.a(new_n11373), .b(new_n11372), .O(new_n11374));
  nor2 g11181(.a(new_n11374), .b(new_n11371), .O(new_n11375));
  nor2 g11182(.a(new_n10892), .b(new_n10885), .O(new_n11376));
  nor2 g11183(.a(new_n11376), .b(new_n11375), .O(new_n11377));
  inv1 g11184(.a(new_n11375), .O(new_n11378));
  inv1 g11185(.a(new_n11376), .O(new_n11379));
  nor2 g11186(.a(new_n11379), .b(new_n11378), .O(new_n11380));
  nor2 g11187(.a(new_n11380), .b(new_n11377), .O(new_n11381));
  inv1 g11188(.a(new_n11381), .O(new_n11382));
  nor2 g11189(.a(new_n10895), .b(new_n194), .O(new_n11383));
  nor2 g11190(.a(new_n11383), .b(new_n10835), .O(new_n11384));
  inv1 g11191(.a(new_n11383), .O(new_n11385));
  nor2 g11192(.a(new_n11385), .b(new_n10836), .O(new_n11386));
  nor2 g11193(.a(new_n11386), .b(new_n11384), .O(new_n11387));
  nor2 g11194(.a(new_n10841), .b(new_n10834), .O(new_n11388));
  nor2 g11195(.a(new_n11388), .b(new_n11387), .O(new_n11389));
  inv1 g11196(.a(new_n11387), .O(new_n11390));
  inv1 g11197(.a(new_n11388), .O(new_n11391));
  nor2 g11198(.a(new_n11391), .b(new_n11390), .O(new_n11392));
  nor2 g11199(.a(new_n11392), .b(new_n11389), .O(new_n11393));
  inv1 g11200(.a(new_n11393), .O(new_n11394));
  nor2 g11201(.a(new_n10853), .b(new_n10846), .O(new_n11395));
  inv1 g11202(.a(new_n11395), .O(new_n11396));
  nor2 g11203(.a(new_n11396), .b(new_n11394), .O(new_n11397));
  nor2 g11204(.a(new_n11395), .b(new_n11393), .O(new_n11398));
  nor2 g11205(.a(new_n11398), .b(new_n11397), .O(new_n11399));
  inv1 g11206(.a(new_n11399), .O(new_n11400));
  nor2 g11207(.a(new_n11400), .b(new_n11382), .O(new_n11401));
  nor2 g11208(.a(new_n11399), .b(new_n11381), .O(new_n11402));
  nor2 g11209(.a(new_n11402), .b(new_n11401), .O(new_n11403));
  inv1 g11210(.a(new_n11403), .O(new_n11404));
  nor2 g11211(.a(new_n11404), .b(new_n11368), .O(new_n11405));
  nor2 g11212(.a(new_n11403), .b(new_n11367), .O(new_n11406));
  nor2 g11213(.a(new_n11406), .b(new_n11405), .O(new_n11407));
  inv1 g11214(.a(new_n11407), .O(new_n11408));
  nor2 g11215(.a(new_n11408), .b(new_n11354), .O(new_n11409));
  nor2 g11216(.a(new_n11407), .b(new_n11353), .O(new_n11410));
  nor2 g11217(.a(new_n11410), .b(new_n11409), .O(new_n11411));
  nor2 g11218(.a(new_n11411), .b(new_n11340), .O(new_n11412));
  inv1 g11219(.a(new_n11411), .O(new_n11413));
  nor2 g11220(.a(new_n11413), .b(new_n11339), .O(new_n11414));
  nor2 g11221(.a(new_n11414), .b(new_n11412), .O(new_n11415));
  inv1 g11222(.a(new_n11415), .O(new_n11416));
  nor2 g11223(.a(new_n10810), .b(new_n10806), .O(new_n11417));
  inv1 g11224(.a(new_n11417), .O(new_n11418));
  nor2 g11225(.a(new_n10975), .b(new_n10970), .O(new_n11419));
  inv1 g11226(.a(new_n11419), .O(new_n11420));
  nor2 g11227(.a(new_n11420), .b(new_n11418), .O(new_n11421));
  nor2 g11228(.a(new_n11419), .b(new_n11417), .O(new_n11422));
  nor2 g11229(.a(new_n11422), .b(new_n11421), .O(new_n11423));
  nor2 g11230(.a(new_n10775), .b(new_n10769), .O(new_n11424));
  inv1 g11231(.a(new_n11424), .O(new_n11425));
  nor2 g11232(.a(new_n11425), .b(new_n11423), .O(new_n11426));
  inv1 g11233(.a(new_n11423), .O(new_n11427));
  nor2 g11234(.a(new_n11424), .b(new_n11427), .O(new_n11428));
  nor2 g11235(.a(new_n11428), .b(new_n11426), .O(new_n11429));
  nor2 g11236(.a(new_n10942), .b(new_n10937), .O(new_n11430));
  inv1 g11237(.a(new_n11430), .O(new_n11431));
  nor2 g11238(.a(new_n11431), .b(new_n11429), .O(new_n11432));
  inv1 g11239(.a(new_n11429), .O(new_n11433));
  nor2 g11240(.a(new_n11430), .b(new_n11433), .O(new_n11434));
  nor2 g11241(.a(new_n11434), .b(new_n11432), .O(new_n11435));
  inv1 g11242(.a(new_n11435), .O(new_n11436));
  nor2 g11243(.a(new_n11436), .b(new_n11416), .O(new_n11437));
  nor2 g11244(.a(new_n11435), .b(new_n11415), .O(new_n11438));
  nor2 g11245(.a(new_n11438), .b(new_n11437), .O(new_n11439));
  inv1 g11246(.a(new_n11439), .O(new_n11440));
  nor2 g11247(.a(new_n11440), .b(new_n11338), .O(new_n11441));
  inv1 g11248(.a(new_n11338), .O(new_n11442));
  nor2 g11249(.a(new_n11439), .b(new_n11442), .O(new_n11443));
  nor2 g11250(.a(new_n11443), .b(new_n11441), .O(new_n11444));
  inv1 g11251(.a(new_n11444), .O(new_n11445));
  nor2 g11252(.a(new_n11445), .b(new_n11337), .O(new_n11446));
  nor2 g11253(.a(new_n11444), .b(new_n11336), .O(new_n11447));
  nor2 g11254(.a(new_n11447), .b(new_n11446), .O(new_n11448));
  inv1 g11255(.a(new_n11448), .O(new_n11449));
  nor2 g11256(.a(new_n11449), .b(new_n11103), .O(new_n11450));
  inv1 g11257(.a(new_n11103), .O(new_n11451));
  nor2 g11258(.a(new_n11448), .b(new_n11451), .O(new_n11452));
  nor2 g11259(.a(new_n11452), .b(new_n11450), .O(new_n11453));
  inv1 g11260(.a(new_n11453), .O(new_n11454));
  nor2 g11261(.a(new_n11098), .b(new_n11094), .O(new_n11455));
  nor2 g11262(.a(new_n11455), .b(new_n11454), .O(new_n11456));
  inv1 g11263(.a(new_n11455), .O(new_n11457));
  nor2 g11264(.a(new_n11457), .b(new_n11453), .O(new_n11458));
  nor2 g11265(.a(new_n11458), .b(new_n11456), .O(new_n11459));
  inv1 g11266(.a(new_n11459), .O(\asquared[63] ));
  nor2 g11267(.a(new_n11446), .b(new_n11441), .O(new_n11461));
  inv1 g11268(.a(new_n11461), .O(new_n11462));
  nor2 g11269(.a(new_n11335), .b(new_n11168), .O(new_n11463));
  inv1 g11270(.a(new_n11463), .O(new_n11464));
  nor2 g11271(.a(new_n11329), .b(new_n11322), .O(new_n11465));
  nor2 g11272(.a(new_n11405), .b(new_n11401), .O(new_n11466));
  inv1 g11273(.a(new_n11466), .O(new_n11467));
  nor2 g11274(.a(new_n11352), .b(new_n11346), .O(new_n11468));
  inv1 g11275(.a(new_n11468), .O(new_n11469));
  nor2 g11276(.a(new_n11469), .b(new_n11467), .O(new_n11470));
  nor2 g11277(.a(new_n11468), .b(new_n11466), .O(new_n11471));
  nor2 g11278(.a(new_n11471), .b(new_n11470), .O(new_n11472));
  nor2 g11279(.a(new_n11139), .b(new_n11133), .O(new_n11473));
  inv1 g11280(.a(new_n11473), .O(new_n11474));
  nor2 g11281(.a(new_n11474), .b(new_n11472), .O(new_n11475));
  inv1 g11282(.a(new_n11472), .O(new_n11476));
  nor2 g11283(.a(new_n11473), .b(new_n11476), .O(new_n11477));
  nor2 g11284(.a(new_n11477), .b(new_n11475), .O(new_n11478));
  inv1 g11285(.a(new_n11478), .O(new_n11479));
  nor2 g11286(.a(new_n11380), .b(new_n11374), .O(new_n11480));
  inv1 g11287(.a(new_n11480), .O(new_n11481));
  nor2 g11288(.a(new_n11125), .b(new_n11110), .O(new_n11482));
  inv1 g11289(.a(new_n11482), .O(new_n11483));
  nor2 g11290(.a(new_n11483), .b(new_n11481), .O(new_n11484));
  nor2 g11291(.a(new_n11482), .b(new_n11480), .O(new_n11485));
  nor2 g11292(.a(new_n11485), .b(new_n11484), .O(new_n11486));
  nor2 g11293(.a(new_n11397), .b(new_n11392), .O(new_n11487));
  inv1 g11294(.a(new_n11487), .O(new_n11488));
  nor2 g11295(.a(new_n11488), .b(new_n11486), .O(new_n11489));
  inv1 g11296(.a(new_n11486), .O(new_n11490));
  nor2 g11297(.a(new_n11487), .b(new_n11490), .O(new_n11491));
  nor2 g11298(.a(new_n11491), .b(new_n11489), .O(new_n11492));
  inv1 g11299(.a(new_n11492), .O(new_n11493));
  nor2 g11300(.a(new_n11318), .b(new_n11264), .O(new_n11494));
  nor2 g11301(.a(new_n11494), .b(new_n11493), .O(new_n11495));
  inv1 g11302(.a(new_n11494), .O(new_n11496));
  nor2 g11303(.a(new_n11496), .b(new_n11492), .O(new_n11497));
  nor2 g11304(.a(new_n11497), .b(new_n11495), .O(new_n11498));
  inv1 g11305(.a(new_n11498), .O(new_n11499));
  nor2 g11306(.a(new_n11279), .b(new_n11272), .O(new_n11500));
  nor2 g11307(.a(new_n11231), .b(new_n11224), .O(new_n11501));
  nor2 g11308(.a(new_n11501), .b(new_n11500), .O(new_n11502));
  inv1 g11309(.a(new_n11500), .O(new_n11503));
  inv1 g11310(.a(new_n11501), .O(new_n11504));
  nor2 g11311(.a(new_n11504), .b(new_n11503), .O(new_n11505));
  nor2 g11312(.a(new_n11505), .b(new_n11502), .O(new_n11506));
  nor2 g11313(.a(new_n11252), .b(new_n11247), .O(new_n11507));
  nor2 g11314(.a(new_n11507), .b(new_n11506), .O(new_n11508));
  inv1 g11315(.a(new_n11506), .O(new_n11509));
  inv1 g11316(.a(new_n11507), .O(new_n11510));
  nor2 g11317(.a(new_n11510), .b(new_n11509), .O(new_n11511));
  nor2 g11318(.a(new_n11511), .b(new_n11508), .O(new_n11512));
  inv1 g11319(.a(new_n11512), .O(new_n11513));
  nor2 g11320(.a(new_n11123), .b(new_n11116), .O(new_n11514));
  nor2 g11321(.a(new_n11208), .b(new_n11200), .O(new_n11515));
  nor2 g11322(.a(new_n11515), .b(new_n11514), .O(new_n11516));
  inv1 g11323(.a(new_n11514), .O(new_n11517));
  inv1 g11324(.a(new_n11515), .O(new_n11518));
  nor2 g11325(.a(new_n11518), .b(new_n11517), .O(new_n11519));
  nor2 g11326(.a(new_n11519), .b(new_n11516), .O(new_n11520));
  nor2 g11327(.a(new_n11195), .b(new_n11189), .O(new_n11521));
  nor2 g11328(.a(new_n11521), .b(new_n11520), .O(new_n11522));
  inv1 g11329(.a(new_n11520), .O(new_n11523));
  inv1 g11330(.a(new_n11521), .O(new_n11524));
  nor2 g11331(.a(new_n11524), .b(new_n11523), .O(new_n11525));
  nor2 g11332(.a(new_n11525), .b(new_n11522), .O(new_n11526));
  nor2 g11333(.a(new_n11366), .b(new_n11360), .O(new_n11527));
  inv1 g11334(.a(new_n11527), .O(new_n11528));
  nor2 g11335(.a(new_n11528), .b(new_n11526), .O(new_n11529));
  inv1 g11336(.a(new_n11526), .O(new_n11530));
  nor2 g11337(.a(new_n11527), .b(new_n11530), .O(new_n11531));
  nor2 g11338(.a(new_n11531), .b(new_n11529), .O(new_n11532));
  inv1 g11339(.a(new_n11532), .O(new_n11533));
  nor2 g11340(.a(new_n11533), .b(new_n11513), .O(new_n11534));
  nor2 g11341(.a(new_n11532), .b(new_n11512), .O(new_n11535));
  nor2 g11342(.a(new_n11535), .b(new_n11534), .O(new_n11536));
  inv1 g11343(.a(new_n11536), .O(new_n11537));
  nor2 g11344(.a(new_n11537), .b(new_n11499), .O(new_n11538));
  nor2 g11345(.a(new_n11536), .b(new_n11498), .O(new_n11539));
  nor2 g11346(.a(new_n11539), .b(new_n11538), .O(new_n11540));
  inv1 g11347(.a(new_n11540), .O(new_n11541));
  nor2 g11348(.a(new_n11541), .b(new_n11479), .O(new_n11542));
  nor2 g11349(.a(new_n11540), .b(new_n11478), .O(new_n11543));
  nor2 g11350(.a(new_n11543), .b(new_n11542), .O(new_n11544));
  inv1 g11351(.a(new_n11544), .O(new_n11545));
  nor2 g11352(.a(new_n11545), .b(new_n11465), .O(new_n11546));
  inv1 g11353(.a(new_n11465), .O(new_n11547));
  nor2 g11354(.a(new_n11544), .b(new_n11547), .O(new_n11548));
  nor2 g11355(.a(new_n11548), .b(new_n11546), .O(new_n11549));
  nor2 g11356(.a(new_n11549), .b(new_n11464), .O(new_n11550));
  inv1 g11357(.a(new_n11549), .O(new_n11551));
  nor2 g11358(.a(new_n11551), .b(new_n11463), .O(new_n11552));
  nor2 g11359(.a(new_n11552), .b(new_n11550), .O(new_n11553));
  nor2 g11360(.a(new_n11437), .b(new_n11434), .O(new_n11554));
  nor2 g11361(.a(new_n11428), .b(new_n11422), .O(new_n11555));
  nor2 g11362(.a(new_n11306), .b(new_n11298), .O(new_n11556));
  nor2 g11363(.a(new_n11182), .b(new_n11177), .O(new_n11557));
  nor2 g11364(.a(new_n11557), .b(new_n11556), .O(new_n11558));
  inv1 g11365(.a(new_n11556), .O(new_n11559));
  inv1 g11366(.a(new_n11557), .O(new_n11560));
  nor2 g11367(.a(new_n11560), .b(new_n11559), .O(new_n11561));
  nor2 g11368(.a(new_n11561), .b(new_n11558), .O(new_n11562));
  nor2 g11369(.a(new_n11291), .b(new_n11284), .O(new_n11563));
  nor2 g11370(.a(new_n11563), .b(new_n11562), .O(new_n11564));
  inv1 g11371(.a(new_n11562), .O(new_n11565));
  inv1 g11372(.a(new_n11563), .O(new_n11566));
  nor2 g11373(.a(new_n11566), .b(new_n11565), .O(new_n11567));
  nor2 g11374(.a(new_n11567), .b(new_n11564), .O(new_n11568));
  nor2 g11375(.a(new_n11315), .b(new_n11308), .O(new_n11569));
  inv1 g11376(.a(new_n11569), .O(new_n11570));
  nor2 g11377(.a(new_n11570), .b(new_n11568), .O(new_n11571));
  inv1 g11378(.a(new_n11568), .O(new_n11572));
  nor2 g11379(.a(new_n11569), .b(new_n11572), .O(new_n11573));
  nor2 g11380(.a(new_n11573), .b(new_n11571), .O(new_n11574));
  nor2 g11381(.a(new_n11261), .b(new_n11254), .O(new_n11575));
  inv1 g11382(.a(new_n11575), .O(new_n11576));
  nor2 g11383(.a(new_n11576), .b(new_n11574), .O(new_n11577));
  inv1 g11384(.a(new_n11574), .O(new_n11578));
  nor2 g11385(.a(new_n11575), .b(new_n11578), .O(new_n11579));
  nor2 g11386(.a(new_n11579), .b(new_n11577), .O(new_n11580));
  nor2 g11387(.a(new_n11155), .b(new_n11149), .O(new_n11581));
  inv1 g11388(.a(new_n11581), .O(new_n11582));
  nor2 g11389(.a(new_n11217), .b(new_n11210), .O(new_n11583));
  inv1 g11390(.a(new_n11583), .O(new_n11584));
  nor2 g11391(.a(new_n11584), .b(new_n11582), .O(new_n11585));
  nor2 g11392(.a(new_n11583), .b(new_n11581), .O(new_n11586));
  nor2 g11393(.a(new_n11586), .b(new_n11585), .O(new_n11587));
  inv1 g11394(.a(new_n11587), .O(new_n11588));
  nor2 g11395(.a(new_n3329), .b(new_n11186), .O(new_n11589));
  nor2 g11396(.a(new_n11589), .b(new_n3057), .O(new_n11590));
  nor2 g11397(.a(\a[32] ), .b(new_n194), .O(new_n11591));
  inv1 g11398(.a(new_n11591), .O(new_n11592));
  nor2 g11399(.a(new_n11592), .b(new_n11186), .O(new_n11593));
  nor2 g11400(.a(new_n11593), .b(new_n11590), .O(new_n11594));
  inv1 g11401(.a(new_n11386), .O(new_n11595));
  inv1 g11402(.a(\a[63] ), .O(new_n11596));
  nor2 g11403(.a(new_n11596), .b(new_n198), .O(new_n11597));
  inv1 g11404(.a(new_n11597), .O(new_n11598));
  nor2 g11405(.a(new_n11598), .b(new_n11595), .O(new_n11599));
  nor2 g11406(.a(new_n11597), .b(new_n11386), .O(new_n11600));
  nor2 g11407(.a(new_n11600), .b(new_n11599), .O(new_n11601));
  inv1 g11408(.a(new_n11601), .O(new_n11602));
  nor2 g11409(.a(new_n11602), .b(new_n11594), .O(new_n11603));
  inv1 g11410(.a(new_n11594), .O(new_n11604));
  nor2 g11411(.a(new_n11601), .b(new_n11604), .O(new_n11605));
  nor2 g11412(.a(new_n11605), .b(new_n11603), .O(new_n11606));
  inv1 g11413(.a(new_n11606), .O(new_n11607));
  nor2 g11414(.a(new_n4366), .b(new_n1903), .O(new_n11608));
  nor2 g11415(.a(new_n11608), .b(new_n11202), .O(new_n11609));
  nor2 g11416(.a(new_n4366), .b(new_n2121), .O(new_n11610));
  inv1 g11417(.a(new_n11610), .O(new_n11611));
  nor2 g11418(.a(new_n11611), .b(new_n10887), .O(new_n11612));
  nor2 g11419(.a(new_n11612), .b(new_n11609), .O(new_n11613));
  inv1 g11420(.a(new_n11613), .O(new_n11614));
  nor2 g11421(.a(new_n11614), .b(new_n11273), .O(new_n11615));
  nor2 g11422(.a(new_n11613), .b(new_n11274), .O(new_n11616));
  nor2 g11423(.a(new_n11616), .b(new_n11615), .O(new_n11617));
  nor2 g11424(.a(new_n3870), .b(new_n2184), .O(new_n11618));
  inv1 g11425(.a(new_n11618), .O(new_n11619));
  nor2 g11426(.a(new_n3722), .b(new_n2433), .O(new_n11620));
  nor2 g11427(.a(new_n11620), .b(new_n11300), .O(new_n11621));
  nor2 g11428(.a(new_n3722), .b(new_n2506), .O(new_n11622));
  inv1 g11429(.a(new_n11622), .O(new_n11623));
  nor2 g11430(.a(new_n11623), .b(new_n11020), .O(new_n11624));
  nor2 g11431(.a(new_n11624), .b(new_n11621), .O(new_n11625));
  nor2 g11432(.a(new_n11625), .b(new_n11619), .O(new_n11626));
  inv1 g11433(.a(new_n11625), .O(new_n11627));
  nor2 g11434(.a(new_n11627), .b(new_n11618), .O(new_n11628));
  nor2 g11435(.a(new_n11628), .b(new_n11626), .O(new_n11629));
  nor2 g11436(.a(new_n11629), .b(new_n11617), .O(new_n11630));
  inv1 g11437(.a(new_n11617), .O(new_n11631));
  inv1 g11438(.a(new_n11629), .O(new_n11632));
  nor2 g11439(.a(new_n11632), .b(new_n11631), .O(new_n11633));
  nor2 g11440(.a(new_n11633), .b(new_n11630), .O(new_n11634));
  inv1 g11441(.a(new_n11634), .O(new_n11635));
  nor2 g11442(.a(new_n11635), .b(new_n11607), .O(new_n11636));
  nor2 g11443(.a(new_n11634), .b(new_n11606), .O(new_n11637));
  nor2 g11444(.a(new_n11637), .b(new_n11636), .O(new_n11638));
  inv1 g11445(.a(new_n11638), .O(new_n11639));
  nor2 g11446(.a(new_n11639), .b(new_n11588), .O(new_n11640));
  nor2 g11447(.a(new_n11638), .b(new_n11587), .O(new_n11641));
  nor2 g11448(.a(new_n11641), .b(new_n11640), .O(new_n11642));
  nor2 g11449(.a(new_n11642), .b(new_n11580), .O(new_n11643));
  inv1 g11450(.a(new_n11580), .O(new_n11644));
  inv1 g11451(.a(new_n11642), .O(new_n11645));
  nor2 g11452(.a(new_n11645), .b(new_n11644), .O(new_n11646));
  nor2 g11453(.a(new_n11646), .b(new_n11643), .O(new_n11647));
  inv1 g11454(.a(new_n11647), .O(new_n11648));
  nor2 g11455(.a(new_n11648), .b(new_n11555), .O(new_n11649));
  inv1 g11456(.a(new_n11555), .O(new_n11650));
  nor2 g11457(.a(new_n11647), .b(new_n11650), .O(new_n11651));
  nor2 g11458(.a(new_n11651), .b(new_n11649), .O(new_n11652));
  inv1 g11459(.a(new_n11652), .O(new_n11653));
  nor2 g11460(.a(new_n11653), .b(new_n11554), .O(new_n11654));
  inv1 g11461(.a(new_n11554), .O(new_n11655));
  nor2 g11462(.a(new_n11652), .b(new_n11655), .O(new_n11656));
  nor2 g11463(.a(new_n11656), .b(new_n11654), .O(new_n11657));
  inv1 g11464(.a(new_n11657), .O(new_n11658));
  nor2 g11465(.a(new_n11414), .b(new_n11409), .O(new_n11659));
  nor2 g11466(.a(new_n11164), .b(new_n11159), .O(new_n11660));
  nor2 g11467(.a(new_n5971), .b(new_n1086), .O(new_n11661));
  nor2 g11468(.a(new_n8476), .b(new_n363), .O(new_n11662));
  nor2 g11469(.a(new_n11662), .b(new_n7285), .O(new_n11663));
  nor2 g11470(.a(new_n8476), .b(new_n941), .O(new_n11664));
  inv1 g11471(.a(new_n11664), .O(new_n11665));
  nor2 g11472(.a(new_n11665), .b(new_n8999), .O(new_n11666));
  nor2 g11473(.a(new_n11666), .b(new_n11663), .O(new_n11667));
  inv1 g11474(.a(new_n11667), .O(new_n11668));
  nor2 g11475(.a(new_n11668), .b(new_n11661), .O(new_n11669));
  inv1 g11476(.a(new_n11661), .O(new_n11670));
  nor2 g11477(.a(new_n11667), .b(new_n11670), .O(new_n11671));
  nor2 g11478(.a(new_n11671), .b(new_n11669), .O(new_n11672));
  nor2 g11479(.a(new_n8170), .b(new_n438), .O(new_n11673));
  inv1 g11480(.a(new_n11673), .O(new_n11674));
  nor2 g11481(.a(new_n6570), .b(new_n847), .O(new_n11675));
  nor2 g11482(.a(new_n8026), .b(new_n502), .O(new_n11676));
  nor2 g11483(.a(new_n11676), .b(new_n11675), .O(new_n11677));
  nor2 g11484(.a(new_n8026), .b(new_n847), .O(new_n11678));
  inv1 g11485(.a(new_n11678), .O(new_n11679));
  nor2 g11486(.a(new_n11679), .b(new_n11236), .O(new_n11680));
  nor2 g11487(.a(new_n11680), .b(new_n11677), .O(new_n11681));
  nor2 g11488(.a(new_n11681), .b(new_n11674), .O(new_n11682));
  inv1 g11489(.a(new_n11681), .O(new_n11683));
  nor2 g11490(.a(new_n11683), .b(new_n11673), .O(new_n11684));
  nor2 g11491(.a(new_n11684), .b(new_n11682), .O(new_n11685));
  nor2 g11492(.a(new_n11685), .b(new_n11672), .O(new_n11686));
  inv1 g11493(.a(new_n11672), .O(new_n11687));
  inv1 g11494(.a(new_n11685), .O(new_n11688));
  nor2 g11495(.a(new_n11688), .b(new_n11687), .O(new_n11689));
  nor2 g11496(.a(new_n11689), .b(new_n11686), .O(new_n11690));
  inv1 g11497(.a(new_n11690), .O(new_n11691));
  nor2 g11498(.a(new_n7537), .b(new_n569), .O(new_n11692));
  nor2 g11499(.a(new_n7294), .b(new_n613), .O(new_n11693));
  nor2 g11500(.a(new_n11693), .b(new_n11692), .O(new_n11694));
  nor2 g11501(.a(new_n7537), .b(new_n613), .O(new_n11695));
  inv1 g11502(.a(new_n11695), .O(new_n11696));
  nor2 g11503(.a(new_n11696), .b(new_n11244), .O(new_n11697));
  nor2 g11504(.a(new_n11697), .b(new_n11694), .O(new_n11698));
  nor2 g11505(.a(new_n11698), .b(new_n9063), .O(new_n11699));
  inv1 g11506(.a(new_n11698), .O(new_n11700));
  nor2 g11507(.a(new_n11700), .b(new_n9062), .O(new_n11701));
  nor2 g11508(.a(new_n11701), .b(new_n11699), .O(new_n11702));
  nor2 g11509(.a(new_n11702), .b(new_n11691), .O(new_n11703));
  inv1 g11510(.a(new_n11702), .O(new_n11704));
  nor2 g11511(.a(new_n11704), .b(new_n11690), .O(new_n11705));
  nor2 g11512(.a(new_n11705), .b(new_n11703), .O(new_n11706));
  inv1 g11513(.a(new_n11706), .O(new_n11707));
  nor2 g11514(.a(new_n5178), .b(new_n1425), .O(new_n11708));
  nor2 g11515(.a(new_n4954), .b(new_n1493), .O(new_n11709));
  nor2 g11516(.a(new_n11709), .b(new_n11708), .O(new_n11710));
  nor2 g11517(.a(new_n5178), .b(new_n1493), .O(new_n11711));
  inv1 g11518(.a(new_n11711), .O(new_n11712));
  nor2 g11519(.a(new_n11712), .b(new_n10915), .O(new_n11713));
  nor2 g11520(.a(new_n11713), .b(new_n11710), .O(new_n11714));
  nor2 g11521(.a(new_n11714), .b(new_n11118), .O(new_n11715));
  inv1 g11522(.a(new_n11714), .O(new_n11716));
  nor2 g11523(.a(new_n11716), .b(new_n11117), .O(new_n11717));
  nor2 g11524(.a(new_n11717), .b(new_n11715), .O(new_n11718));
  nor2 g11525(.a(new_n10895), .b(new_n196), .O(new_n11719));
  inv1 g11526(.a(new_n11719), .O(new_n11720));
  nor2 g11527(.a(new_n10468), .b(new_n203), .O(new_n11721));
  nor2 g11528(.a(new_n10320), .b(new_n214), .O(new_n11722));
  nor2 g11529(.a(new_n11722), .b(new_n11721), .O(new_n11723));
  nor2 g11530(.a(new_n10468), .b(new_n214), .O(new_n11724));
  inv1 g11531(.a(new_n11724), .O(new_n11725));
  nor2 g11532(.a(new_n11725), .b(new_n11114), .O(new_n11726));
  nor2 g11533(.a(new_n11726), .b(new_n11723), .O(new_n11727));
  nor2 g11534(.a(new_n11727), .b(new_n11720), .O(new_n11728));
  inv1 g11535(.a(new_n11727), .O(new_n11729));
  nor2 g11536(.a(new_n11729), .b(new_n11719), .O(new_n11730));
  nor2 g11537(.a(new_n11730), .b(new_n11728), .O(new_n11731));
  nor2 g11538(.a(new_n11240), .b(new_n11235), .O(new_n11732));
  inv1 g11539(.a(new_n11732), .O(new_n11733));
  nor2 g11540(.a(new_n11733), .b(new_n11731), .O(new_n11734));
  inv1 g11541(.a(new_n11731), .O(new_n11735));
  nor2 g11542(.a(new_n11732), .b(new_n11735), .O(new_n11736));
  nor2 g11543(.a(new_n11736), .b(new_n11734), .O(new_n11737));
  inv1 g11544(.a(new_n11737), .O(new_n11738));
  nor2 g11545(.a(new_n11738), .b(new_n11718), .O(new_n11739));
  inv1 g11546(.a(new_n11718), .O(new_n11740));
  nor2 g11547(.a(new_n11737), .b(new_n11740), .O(new_n11741));
  nor2 g11548(.a(new_n11741), .b(new_n11739), .O(new_n11742));
  inv1 g11549(.a(new_n11742), .O(new_n11743));
  nor2 g11550(.a(new_n8946), .b(new_n322), .O(new_n11744));
  nor2 g11551(.a(new_n5796), .b(new_n1199), .O(new_n11745));
  nor2 g11552(.a(new_n11745), .b(new_n11744), .O(new_n11746));
  nor2 g11553(.a(new_n8946), .b(new_n1199), .O(new_n11747));
  inv1 g11554(.a(new_n11747), .O(new_n11748));
  nor2 g11555(.a(new_n11748), .b(new_n11285), .O(new_n11749));
  nor2 g11556(.a(new_n11749), .b(new_n11746), .O(new_n11750));
  nor2 g11557(.a(new_n11750), .b(new_n11226), .O(new_n11751));
  inv1 g11558(.a(new_n11750), .O(new_n11752));
  nor2 g11559(.a(new_n11752), .b(new_n11225), .O(new_n11753));
  nor2 g11560(.a(new_n11753), .b(new_n11751), .O(new_n11754));
  nor2 g11561(.a(new_n3057), .b(new_n2826), .O(new_n11755));
  nor2 g11562(.a(new_n3231), .b(new_n2660), .O(new_n11756));
  nor2 g11563(.a(new_n11756), .b(new_n11755), .O(new_n11757));
  inv1 g11564(.a(new_n11755), .O(new_n11758));
  inv1 g11565(.a(new_n11756), .O(new_n11759));
  nor2 g11566(.a(new_n11759), .b(new_n11758), .O(new_n11760));
  nor2 g11567(.a(new_n11760), .b(new_n11757), .O(new_n11761));
  nor2 g11568(.a(new_n11761), .b(new_n10848), .O(new_n11762));
  inv1 g11569(.a(new_n11761), .O(new_n11763));
  nor2 g11570(.a(new_n11763), .b(new_n10847), .O(new_n11764));
  nor2 g11571(.a(new_n11764), .b(new_n11762), .O(new_n11765));
  nor2 g11572(.a(new_n4682), .b(new_n1647), .O(new_n11766));
  inv1 g11573(.a(new_n11766), .O(new_n11767));
  nor2 g11574(.a(new_n9658), .b(new_n257), .O(new_n11768));
  nor2 g11575(.a(new_n5393), .b(new_n1297), .O(new_n11769));
  nor2 g11576(.a(new_n11769), .b(new_n11768), .O(new_n11770));
  inv1 g11577(.a(new_n11768), .O(new_n11771));
  inv1 g11578(.a(new_n11769), .O(new_n11772));
  nor2 g11579(.a(new_n11772), .b(new_n11771), .O(new_n11773));
  nor2 g11580(.a(new_n11773), .b(new_n11770), .O(new_n11774));
  inv1 g11581(.a(new_n11774), .O(new_n11775));
  nor2 g11582(.a(new_n11775), .b(new_n11767), .O(new_n11776));
  nor2 g11583(.a(new_n11774), .b(new_n11766), .O(new_n11777));
  nor2 g11584(.a(new_n11777), .b(new_n11776), .O(new_n11778));
  inv1 g11585(.a(new_n11778), .O(new_n11779));
  nor2 g11586(.a(new_n11779), .b(new_n11765), .O(new_n11780));
  inv1 g11587(.a(new_n11765), .O(new_n11781));
  nor2 g11588(.a(new_n11778), .b(new_n11781), .O(new_n11782));
  nor2 g11589(.a(new_n11782), .b(new_n11780), .O(new_n11783));
  inv1 g11590(.a(new_n11783), .O(new_n11784));
  nor2 g11591(.a(new_n11784), .b(new_n11754), .O(new_n11785));
  inv1 g11592(.a(new_n11754), .O(new_n11786));
  nor2 g11593(.a(new_n11783), .b(new_n11786), .O(new_n11787));
  nor2 g11594(.a(new_n11787), .b(new_n11785), .O(new_n11788));
  inv1 g11595(.a(new_n11788), .O(new_n11789));
  nor2 g11596(.a(new_n11789), .b(new_n11743), .O(new_n11790));
  nor2 g11597(.a(new_n11788), .b(new_n11742), .O(new_n11791));
  nor2 g11598(.a(new_n11791), .b(new_n11790), .O(new_n11792));
  inv1 g11599(.a(new_n11792), .O(new_n11793));
  nor2 g11600(.a(new_n11793), .b(new_n11707), .O(new_n11794));
  nor2 g11601(.a(new_n11792), .b(new_n11706), .O(new_n11795));
  nor2 g11602(.a(new_n11795), .b(new_n11794), .O(new_n11796));
  inv1 g11603(.a(new_n11796), .O(new_n11797));
  nor2 g11604(.a(new_n11797), .b(new_n11660), .O(new_n11798));
  inv1 g11605(.a(new_n11660), .O(new_n11799));
  nor2 g11606(.a(new_n11796), .b(new_n11799), .O(new_n11800));
  nor2 g11607(.a(new_n11800), .b(new_n11798), .O(new_n11801));
  inv1 g11608(.a(new_n11801), .O(new_n11802));
  nor2 g11609(.a(new_n11802), .b(new_n11659), .O(new_n11803));
  inv1 g11610(.a(new_n11659), .O(new_n11804));
  nor2 g11611(.a(new_n11801), .b(new_n11804), .O(new_n11805));
  nor2 g11612(.a(new_n11805), .b(new_n11803), .O(new_n11806));
  inv1 g11613(.a(new_n11806), .O(new_n11807));
  nor2 g11614(.a(new_n11807), .b(new_n11658), .O(new_n11808));
  nor2 g11615(.a(new_n11806), .b(new_n11657), .O(new_n11809));
  nor2 g11616(.a(new_n11809), .b(new_n11808), .O(new_n11810));
  nor2 g11617(.a(new_n11810), .b(new_n11553), .O(new_n11811));
  inv1 g11618(.a(new_n11553), .O(new_n11812));
  inv1 g11619(.a(new_n11810), .O(new_n11813));
  nor2 g11620(.a(new_n11813), .b(new_n11812), .O(new_n11814));
  nor2 g11621(.a(new_n11814), .b(new_n11811), .O(new_n11815));
  nor2 g11622(.a(new_n11815), .b(new_n11462), .O(new_n11816));
  inv1 g11623(.a(new_n11815), .O(new_n11817));
  nor2 g11624(.a(new_n11817), .b(new_n11461), .O(new_n11818));
  nor2 g11625(.a(new_n11818), .b(new_n11816), .O(new_n11819));
  inv1 g11626(.a(new_n11819), .O(new_n11820));
  nor2 g11627(.a(new_n11456), .b(new_n11452), .O(new_n11821));
  nor2 g11628(.a(new_n11821), .b(new_n11820), .O(new_n11822));
  inv1 g11629(.a(new_n11821), .O(new_n11823));
  nor2 g11630(.a(new_n11823), .b(new_n11819), .O(new_n11824));
  nor2 g11631(.a(new_n11824), .b(new_n11822), .O(new_n11825));
  inv1 g11632(.a(new_n11825), .O(\asquared[64] ));
  nor2 g11633(.a(new_n11546), .b(new_n11542), .O(new_n11827));
  nor2 g11634(.a(new_n11701), .b(new_n11694), .O(new_n11828));
  nor2 g11635(.a(new_n11615), .b(new_n11609), .O(new_n11829));
  nor2 g11636(.a(new_n11829), .b(new_n11828), .O(new_n11830));
  inv1 g11637(.a(new_n11828), .O(new_n11831));
  inv1 g11638(.a(new_n11829), .O(new_n11832));
  nor2 g11639(.a(new_n11832), .b(new_n11831), .O(new_n11833));
  nor2 g11640(.a(new_n11833), .b(new_n11830), .O(new_n11834));
  nor2 g11641(.a(new_n11684), .b(new_n11677), .O(new_n11835));
  nor2 g11642(.a(new_n11835), .b(new_n11834), .O(new_n11836));
  inv1 g11643(.a(new_n11834), .O(new_n11837));
  inv1 g11644(.a(new_n11835), .O(new_n11838));
  nor2 g11645(.a(new_n11838), .b(new_n11837), .O(new_n11839));
  nor2 g11646(.a(new_n11839), .b(new_n11836), .O(new_n11840));
  nor2 g11647(.a(new_n11785), .b(new_n11780), .O(new_n11841));
  inv1 g11648(.a(new_n11841), .O(new_n11842));
  nor2 g11649(.a(new_n11842), .b(new_n11840), .O(new_n11843));
  inv1 g11650(.a(new_n11840), .O(new_n11844));
  nor2 g11651(.a(new_n11841), .b(new_n11844), .O(new_n11845));
  nor2 g11652(.a(new_n11845), .b(new_n11843), .O(new_n11846));
  nor2 g11653(.a(new_n11703), .b(new_n11686), .O(new_n11847));
  inv1 g11654(.a(new_n11847), .O(new_n11848));
  nor2 g11655(.a(new_n11848), .b(new_n11846), .O(new_n11849));
  inv1 g11656(.a(new_n11846), .O(new_n11850));
  nor2 g11657(.a(new_n11847), .b(new_n11850), .O(new_n11851));
  nor2 g11658(.a(new_n11851), .b(new_n11849), .O(new_n11852));
  nor2 g11659(.a(new_n11477), .b(new_n11471), .O(new_n11853));
  inv1 g11660(.a(new_n11853), .O(new_n11854));
  nor2 g11661(.a(new_n11854), .b(new_n11852), .O(new_n11855));
  inv1 g11662(.a(new_n11852), .O(new_n11856));
  nor2 g11663(.a(new_n11853), .b(new_n11856), .O(new_n11857));
  nor2 g11664(.a(new_n11857), .b(new_n11855), .O(new_n11858));
  nor2 g11665(.a(new_n11491), .b(new_n11485), .O(new_n11859));
  inv1 g11666(.a(new_n11859), .O(new_n11860));
  nor2 g11667(.a(new_n11739), .b(new_n11734), .O(new_n11861));
  inv1 g11668(.a(new_n11861), .O(new_n11862));
  nor2 g11669(.a(new_n11862), .b(new_n11860), .O(new_n11863));
  nor2 g11670(.a(new_n11861), .b(new_n11859), .O(new_n11864));
  nor2 g11671(.a(new_n11864), .b(new_n11863), .O(new_n11865));
  inv1 g11672(.a(new_n11865), .O(new_n11866));
  nor2 g11673(.a(new_n11764), .b(new_n11757), .O(new_n11867));
  inv1 g11674(.a(new_n11867), .O(new_n11868));
  inv1 g11675(.a(new_n11589), .O(new_n11869));
  nor2 g11676(.a(new_n11869), .b(new_n11596), .O(new_n11870));
  nor2 g11677(.a(new_n11186), .b(new_n3057), .O(new_n11871));
  nor2 g11678(.a(new_n11871), .b(\a[63] ), .O(new_n11872));
  nor2 g11679(.a(new_n11872), .b(new_n194), .O(new_n11873));
  inv1 g11680(.a(new_n11873), .O(new_n11874));
  nor2 g11681(.a(new_n11874), .b(new_n11870), .O(new_n11875));
  inv1 g11682(.a(new_n11875), .O(new_n11876));
  nor2 g11683(.a(new_n11876), .b(new_n11868), .O(new_n11877));
  nor2 g11684(.a(new_n11875), .b(new_n11867), .O(new_n11878));
  nor2 g11685(.a(new_n11878), .b(new_n11877), .O(new_n11879));
  inv1 g11686(.a(new_n11879), .O(new_n11880));
  nor2 g11687(.a(new_n8170), .b(new_n502), .O(new_n11881));
  nor2 g11688(.a(new_n8026), .b(new_n569), .O(new_n11882));
  nor2 g11689(.a(new_n11882), .b(new_n11881), .O(new_n11883));
  inv1 g11690(.a(new_n11676), .O(new_n11884));
  nor2 g11691(.a(new_n8170), .b(new_n569), .O(new_n11885));
  inv1 g11692(.a(new_n11885), .O(new_n11886));
  nor2 g11693(.a(new_n11886), .b(new_n11884), .O(new_n11887));
  nor2 g11694(.a(new_n11887), .b(new_n11883), .O(new_n11888));
  nor2 g11695(.a(new_n11888), .b(new_n11696), .O(new_n11889));
  inv1 g11696(.a(new_n11888), .O(new_n11890));
  nor2 g11697(.a(new_n11890), .b(new_n11695), .O(new_n11891));
  nor2 g11698(.a(new_n11891), .b(new_n11889), .O(new_n11892));
  nor2 g11699(.a(new_n8946), .b(new_n363), .O(new_n11893));
  inv1 g11700(.a(new_n11893), .O(new_n11894));
  nor2 g11701(.a(new_n8476), .b(new_n438), .O(new_n11895));
  nor2 g11702(.a(new_n11895), .b(new_n10294), .O(new_n11896));
  inv1 g11703(.a(new_n11895), .O(new_n11897));
  nor2 g11704(.a(new_n11897), .b(new_n10295), .O(new_n11898));
  nor2 g11705(.a(new_n11898), .b(new_n11896), .O(new_n11899));
  nor2 g11706(.a(new_n11899), .b(new_n11894), .O(new_n11900));
  inv1 g11707(.a(new_n11899), .O(new_n11901));
  nor2 g11708(.a(new_n11901), .b(new_n11893), .O(new_n11902));
  nor2 g11709(.a(new_n11902), .b(new_n11900), .O(new_n11903));
  nor2 g11710(.a(new_n11903), .b(new_n11892), .O(new_n11904));
  inv1 g11711(.a(new_n11892), .O(new_n11905));
  inv1 g11712(.a(new_n11903), .O(new_n11906));
  nor2 g11713(.a(new_n11906), .b(new_n11905), .O(new_n11907));
  nor2 g11714(.a(new_n11907), .b(new_n11904), .O(new_n11908));
  inv1 g11715(.a(new_n11908), .O(new_n11909));
  nor2 g11716(.a(new_n11909), .b(new_n11880), .O(new_n11910));
  nor2 g11717(.a(new_n11908), .b(new_n11879), .O(new_n11911));
  nor2 g11718(.a(new_n11911), .b(new_n11910), .O(new_n11912));
  inv1 g11719(.a(new_n11912), .O(new_n11913));
  nor2 g11720(.a(new_n11913), .b(new_n11866), .O(new_n11914));
  nor2 g11721(.a(new_n11912), .b(new_n11865), .O(new_n11915));
  nor2 g11722(.a(new_n11915), .b(new_n11914), .O(new_n11916));
  nor2 g11723(.a(new_n11916), .b(new_n11858), .O(new_n11917));
  inv1 g11724(.a(new_n11858), .O(new_n11918));
  inv1 g11725(.a(new_n11916), .O(new_n11919));
  nor2 g11726(.a(new_n11919), .b(new_n11918), .O(new_n11920));
  nor2 g11727(.a(new_n11920), .b(new_n11917), .O(new_n11921));
  inv1 g11728(.a(new_n11921), .O(new_n11922));
  nor2 g11729(.a(new_n11922), .b(new_n11827), .O(new_n11923));
  inv1 g11730(.a(new_n11827), .O(new_n11924));
  nor2 g11731(.a(new_n11921), .b(new_n11924), .O(new_n11925));
  nor2 g11732(.a(new_n11925), .b(new_n11923), .O(new_n11926));
  inv1 g11733(.a(new_n11926), .O(new_n11927));
  nor2 g11734(.a(new_n11538), .b(new_n11495), .O(new_n11928));
  nor2 g11735(.a(new_n10895), .b(new_n203), .O(new_n11929));
  nor2 g11736(.a(new_n11929), .b(new_n11724), .O(new_n11930));
  inv1 g11737(.a(new_n11721), .O(new_n11931));
  nor2 g11738(.a(new_n10895), .b(new_n214), .O(new_n11932));
  inv1 g11739(.a(new_n11932), .O(new_n11933));
  nor2 g11740(.a(new_n11933), .b(new_n11931), .O(new_n11934));
  nor2 g11741(.a(new_n11934), .b(new_n11930), .O(new_n11935));
  nor2 g11742(.a(new_n11935), .b(new_n11191), .O(new_n11936));
  inv1 g11743(.a(new_n11935), .O(new_n11937));
  nor2 g11744(.a(new_n11937), .b(new_n11190), .O(new_n11938));
  nor2 g11745(.a(new_n11938), .b(new_n11936), .O(new_n11939));
  nor2 g11746(.a(new_n6274), .b(new_n1086), .O(new_n11940));
  nor2 g11747(.a(new_n5971), .b(new_n1199), .O(new_n11941));
  nor2 g11748(.a(new_n11941), .b(new_n11940), .O(new_n11942));
  nor2 g11749(.a(new_n6274), .b(new_n1199), .O(new_n11943));
  inv1 g11750(.a(new_n11943), .O(new_n11944));
  nor2 g11751(.a(new_n11944), .b(new_n11670), .O(new_n11945));
  nor2 g11752(.a(new_n11945), .b(new_n11942), .O(new_n11946));
  nor2 g11753(.a(new_n11946), .b(new_n10901), .O(new_n11947));
  inv1 g11754(.a(new_n11946), .O(new_n11948));
  nor2 g11755(.a(new_n11948), .b(new_n10900), .O(new_n11949));
  nor2 g11756(.a(new_n11949), .b(new_n11947), .O(new_n11950));
  nor2 g11757(.a(new_n11603), .b(new_n11599), .O(new_n11951));
  nor2 g11758(.a(new_n11951), .b(new_n11950), .O(new_n11952));
  inv1 g11759(.a(new_n11950), .O(new_n11953));
  inv1 g11760(.a(new_n11951), .O(new_n11954));
  nor2 g11761(.a(new_n11954), .b(new_n11953), .O(new_n11955));
  nor2 g11762(.a(new_n11955), .b(new_n11952), .O(new_n11956));
  inv1 g11763(.a(new_n11956), .O(new_n11957));
  nor2 g11764(.a(new_n11957), .b(new_n11939), .O(new_n11958));
  inv1 g11765(.a(new_n11939), .O(new_n11959));
  nor2 g11766(.a(new_n11956), .b(new_n11959), .O(new_n11960));
  nor2 g11767(.a(new_n11960), .b(new_n11958), .O(new_n11961));
  inv1 g11768(.a(new_n11961), .O(new_n11962));
  nor2 g11769(.a(new_n7294), .b(new_n699), .O(new_n11963));
  inv1 g11770(.a(new_n11963), .O(new_n11964));
  nor2 g11771(.a(new_n3231), .b(new_n2826), .O(new_n11965));
  nor2 g11772(.a(new_n3533), .b(new_n2660), .O(new_n11966));
  nor2 g11773(.a(new_n11966), .b(new_n11965), .O(new_n11967));
  nor2 g11774(.a(new_n3533), .b(new_n2826), .O(new_n11968));
  inv1 g11775(.a(new_n11968), .O(new_n11969));
  nor2 g11776(.a(new_n11969), .b(new_n11759), .O(new_n11970));
  nor2 g11777(.a(new_n11970), .b(new_n11967), .O(new_n11971));
  nor2 g11778(.a(new_n11971), .b(new_n11964), .O(new_n11972));
  inv1 g11779(.a(new_n11971), .O(new_n11973));
  nor2 g11780(.a(new_n11973), .b(new_n11963), .O(new_n11974));
  nor2 g11781(.a(new_n11974), .b(new_n11972), .O(new_n11975));
  inv1 g11782(.a(new_n11975), .O(new_n11976));
  nor2 g11783(.a(new_n9156), .b(new_n322), .O(new_n11977));
  nor2 g11784(.a(new_n11977), .b(new_n8176), .O(new_n11978));
  nor2 g11785(.a(new_n9156), .b(new_n847), .O(new_n11979));
  inv1 g11786(.a(new_n11979), .O(new_n11980));
  nor2 g11787(.a(new_n11980), .b(new_n8868), .O(new_n11981));
  nor2 g11788(.a(new_n11981), .b(new_n11978), .O(new_n11982));
  inv1 g11789(.a(new_n11982), .O(new_n11983));
  nor2 g11790(.a(new_n11983), .b(new_n11610), .O(new_n11984));
  nor2 g11791(.a(new_n11982), .b(new_n11611), .O(new_n11985));
  nor2 g11792(.a(new_n11985), .b(new_n11984), .O(new_n11986));
  nor2 g11793(.a(new_n4093), .b(new_n2184), .O(new_n11987));
  inv1 g11794(.a(new_n11987), .O(new_n11988));
  nor2 g11795(.a(new_n3870), .b(new_n2433), .O(new_n11989));
  nor2 g11796(.a(new_n11989), .b(new_n11622), .O(new_n11990));
  inv1 g11797(.a(new_n11620), .O(new_n11991));
  nor2 g11798(.a(new_n3870), .b(new_n2506), .O(new_n11992));
  inv1 g11799(.a(new_n11992), .O(new_n11993));
  nor2 g11800(.a(new_n11993), .b(new_n11991), .O(new_n11994));
  nor2 g11801(.a(new_n11994), .b(new_n11990), .O(new_n11995));
  nor2 g11802(.a(new_n11995), .b(new_n11988), .O(new_n11996));
  inv1 g11803(.a(new_n11995), .O(new_n11997));
  nor2 g11804(.a(new_n11997), .b(new_n11987), .O(new_n11998));
  nor2 g11805(.a(new_n11998), .b(new_n11996), .O(new_n11999));
  nor2 g11806(.a(new_n11999), .b(new_n11986), .O(new_n12000));
  inv1 g11807(.a(new_n11986), .O(new_n12001));
  inv1 g11808(.a(new_n11999), .O(new_n12002));
  nor2 g11809(.a(new_n12002), .b(new_n12001), .O(new_n12003));
  nor2 g11810(.a(new_n12003), .b(new_n12000), .O(new_n12004));
  nor2 g11811(.a(new_n12004), .b(new_n11976), .O(new_n12005));
  inv1 g11812(.a(new_n12004), .O(new_n12006));
  nor2 g11813(.a(new_n12006), .b(new_n11975), .O(new_n12007));
  nor2 g11814(.a(new_n12007), .b(new_n12005), .O(new_n12008));
  inv1 g11815(.a(new_n12008), .O(new_n12009));
  nor2 g11816(.a(new_n12009), .b(new_n11962), .O(new_n12010));
  nor2 g11817(.a(new_n12008), .b(new_n11961), .O(new_n12011));
  nor2 g11818(.a(new_n12011), .b(new_n12010), .O(new_n12012));
  inv1 g11819(.a(new_n12012), .O(new_n12013));
  nor2 g11820(.a(new_n4954), .b(new_n1647), .O(new_n12014));
  inv1 g11821(.a(new_n12014), .O(new_n12015));
  nor2 g11822(.a(new_n4682), .b(new_n1736), .O(new_n12016));
  nor2 g11823(.a(new_n4425), .b(new_n1903), .O(new_n12017));
  nor2 g11824(.a(new_n12017), .b(new_n12016), .O(new_n12018));
  nor2 g11825(.a(new_n4682), .b(new_n1903), .O(new_n12019));
  inv1 g11826(.a(new_n12019), .O(new_n12020));
  nor2 g11827(.a(new_n12020), .b(new_n11274), .O(new_n12021));
  nor2 g11828(.a(new_n12021), .b(new_n12018), .O(new_n12022));
  nor2 g11829(.a(new_n12022), .b(new_n12015), .O(new_n12023));
  inv1 g11830(.a(new_n12022), .O(new_n12024));
  nor2 g11831(.a(new_n12024), .b(new_n12014), .O(new_n12025));
  nor2 g11832(.a(new_n12025), .b(new_n12023), .O(new_n12026));
  inv1 g11833(.a(new_n12026), .O(new_n12027));
  nor2 g11834(.a(new_n9873), .b(new_n257), .O(new_n12028));
  nor2 g11835(.a(new_n6570), .b(new_n941), .O(new_n12029));
  nor2 g11836(.a(new_n9658), .b(new_n295), .O(new_n12030));
  nor2 g11837(.a(new_n12030), .b(new_n12029), .O(new_n12031));
  nor2 g11838(.a(new_n9658), .b(new_n941), .O(new_n12032));
  inv1 g11839(.a(new_n12032), .O(new_n12033));
  nor2 g11840(.a(new_n12033), .b(new_n8638), .O(new_n12034));
  nor2 g11841(.a(new_n12034), .b(new_n12031), .O(new_n12035));
  inv1 g11842(.a(new_n12035), .O(new_n12036));
  nor2 g11843(.a(new_n12036), .b(new_n12028), .O(new_n12037));
  inv1 g11844(.a(new_n12028), .O(new_n12038));
  nor2 g11845(.a(new_n12035), .b(new_n12038), .O(new_n12039));
  nor2 g11846(.a(new_n12039), .b(new_n12037), .O(new_n12040));
  nor2 g11847(.a(new_n5796), .b(new_n1297), .O(new_n12041));
  inv1 g11848(.a(new_n12041), .O(new_n12042));
  nor2 g11849(.a(new_n5393), .b(new_n1425), .O(new_n12043));
  nor2 g11850(.a(new_n12043), .b(new_n11711), .O(new_n12044));
  inv1 g11851(.a(new_n11708), .O(new_n12045));
  nor2 g11852(.a(new_n5393), .b(new_n1493), .O(new_n12046));
  inv1 g11853(.a(new_n12046), .O(new_n12047));
  nor2 g11854(.a(new_n12047), .b(new_n12045), .O(new_n12048));
  nor2 g11855(.a(new_n12048), .b(new_n12044), .O(new_n12049));
  nor2 g11856(.a(new_n12049), .b(new_n12042), .O(new_n12050));
  inv1 g11857(.a(new_n12049), .O(new_n12051));
  nor2 g11858(.a(new_n12051), .b(new_n12041), .O(new_n12052));
  nor2 g11859(.a(new_n12052), .b(new_n12050), .O(new_n12053));
  nor2 g11860(.a(new_n12053), .b(new_n12040), .O(new_n12054));
  inv1 g11861(.a(new_n12040), .O(new_n12055));
  inv1 g11862(.a(new_n12053), .O(new_n12056));
  nor2 g11863(.a(new_n12056), .b(new_n12055), .O(new_n12057));
  nor2 g11864(.a(new_n12057), .b(new_n12054), .O(new_n12058));
  nor2 g11865(.a(new_n12058), .b(new_n12027), .O(new_n12059));
  inv1 g11866(.a(new_n12058), .O(new_n12060));
  nor2 g11867(.a(new_n12060), .b(new_n12026), .O(new_n12061));
  nor2 g11868(.a(new_n12061), .b(new_n12059), .O(new_n12062));
  inv1 g11869(.a(new_n12062), .O(new_n12063));
  nor2 g11870(.a(new_n12063), .b(new_n12013), .O(new_n12064));
  nor2 g11871(.a(new_n12062), .b(new_n12012), .O(new_n12065));
  nor2 g11872(.a(new_n12065), .b(new_n12064), .O(new_n12066));
  inv1 g11873(.a(new_n12066), .O(new_n12067));
  nor2 g11874(.a(new_n12067), .b(new_n11928), .O(new_n12068));
  inv1 g11875(.a(new_n11928), .O(new_n12069));
  nor2 g11876(.a(new_n12066), .b(new_n12069), .O(new_n12070));
  nor2 g11877(.a(new_n12070), .b(new_n12068), .O(new_n12071));
  inv1 g11878(.a(new_n12071), .O(new_n12072));
  nor2 g11879(.a(new_n11511), .b(new_n11505), .O(new_n12073));
  inv1 g11880(.a(new_n12073), .O(new_n12074));
  nor2 g11881(.a(new_n11567), .b(new_n11561), .O(new_n12075));
  inv1 g11882(.a(new_n12075), .O(new_n12076));
  nor2 g11883(.a(new_n12076), .b(new_n12074), .O(new_n12077));
  nor2 g11884(.a(new_n12075), .b(new_n12073), .O(new_n12078));
  nor2 g11885(.a(new_n12078), .b(new_n12077), .O(new_n12079));
  nor2 g11886(.a(new_n11525), .b(new_n11519), .O(new_n12080));
  inv1 g11887(.a(new_n12080), .O(new_n12081));
  nor2 g11888(.a(new_n12081), .b(new_n12079), .O(new_n12082));
  inv1 g11889(.a(new_n12079), .O(new_n12083));
  nor2 g11890(.a(new_n12080), .b(new_n12083), .O(new_n12084));
  nor2 g11891(.a(new_n12084), .b(new_n12082), .O(new_n12085));
  inv1 g11892(.a(new_n12085), .O(new_n12086));
  nor2 g11893(.a(new_n11579), .b(new_n11573), .O(new_n12087));
  nor2 g11894(.a(new_n11534), .b(new_n11531), .O(new_n12088));
  nor2 g11895(.a(new_n12088), .b(new_n12087), .O(new_n12089));
  inv1 g11896(.a(new_n12087), .O(new_n12090));
  inv1 g11897(.a(new_n12088), .O(new_n12091));
  nor2 g11898(.a(new_n12091), .b(new_n12090), .O(new_n12092));
  nor2 g11899(.a(new_n12092), .b(new_n12089), .O(new_n12093));
  inv1 g11900(.a(new_n12093), .O(new_n12094));
  nor2 g11901(.a(new_n12094), .b(new_n12086), .O(new_n12095));
  nor2 g11902(.a(new_n12093), .b(new_n12085), .O(new_n12096));
  nor2 g11903(.a(new_n12096), .b(new_n12095), .O(new_n12097));
  inv1 g11904(.a(new_n12097), .O(new_n12098));
  nor2 g11905(.a(new_n12098), .b(new_n12072), .O(new_n12099));
  nor2 g11906(.a(new_n12097), .b(new_n12071), .O(new_n12100));
  nor2 g11907(.a(new_n12100), .b(new_n12099), .O(new_n12101));
  inv1 g11908(.a(new_n12101), .O(new_n12102));
  nor2 g11909(.a(new_n12102), .b(new_n11927), .O(new_n12103));
  nor2 g11910(.a(new_n12101), .b(new_n11926), .O(new_n12104));
  nor2 g11911(.a(new_n12104), .b(new_n12103), .O(new_n12105));
  inv1 g11912(.a(new_n12105), .O(new_n12106));
  nor2 g11913(.a(new_n11808), .b(new_n11654), .O(new_n12107));
  nor2 g11914(.a(new_n11803), .b(new_n11798), .O(new_n12108));
  nor2 g11915(.a(new_n11649), .b(new_n11646), .O(new_n12109));
  nor2 g11916(.a(new_n11794), .b(new_n11790), .O(new_n12110));
  inv1 g11917(.a(new_n12110), .O(new_n12111));
  nor2 g11918(.a(new_n11640), .b(new_n11586), .O(new_n12112));
  inv1 g11919(.a(new_n12112), .O(new_n12113));
  nor2 g11920(.a(new_n12113), .b(new_n12111), .O(new_n12114));
  nor2 g11921(.a(new_n12112), .b(new_n12110), .O(new_n12115));
  nor2 g11922(.a(new_n12115), .b(new_n12114), .O(new_n12116));
  nor2 g11923(.a(new_n11636), .b(new_n11630), .O(new_n12117));
  nor2 g11924(.a(new_n11776), .b(new_n11773), .O(new_n12118));
  inv1 g11925(.a(new_n12118), .O(new_n12119));
  nor2 g11926(.a(new_n11669), .b(new_n11663), .O(new_n12120));
  nor2 g11927(.a(new_n12120), .b(new_n12119), .O(new_n12121));
  inv1 g11928(.a(new_n12120), .O(new_n12122));
  nor2 g11929(.a(new_n12122), .b(new_n12118), .O(new_n12123));
  nor2 g11930(.a(new_n12123), .b(new_n12121), .O(new_n12124));
  nor2 g11931(.a(new_n11628), .b(new_n11621), .O(new_n12125));
  nor2 g11932(.a(new_n12125), .b(new_n12124), .O(new_n12126));
  inv1 g11933(.a(new_n12124), .O(new_n12127));
  inv1 g11934(.a(new_n12125), .O(new_n12128));
  nor2 g11935(.a(new_n12128), .b(new_n12127), .O(new_n12129));
  nor2 g11936(.a(new_n12129), .b(new_n12126), .O(new_n12130));
  nor2 g11937(.a(new_n11730), .b(new_n11723), .O(new_n12131));
  nor2 g11938(.a(new_n11717), .b(new_n11710), .O(new_n12132));
  nor2 g11939(.a(new_n12132), .b(new_n12131), .O(new_n12133));
  inv1 g11940(.a(new_n12131), .O(new_n12134));
  inv1 g11941(.a(new_n12132), .O(new_n12135));
  nor2 g11942(.a(new_n12135), .b(new_n12134), .O(new_n12136));
  nor2 g11943(.a(new_n12136), .b(new_n12133), .O(new_n12137));
  nor2 g11944(.a(new_n11753), .b(new_n11746), .O(new_n12138));
  nor2 g11945(.a(new_n12138), .b(new_n12137), .O(new_n12139));
  inv1 g11946(.a(new_n12137), .O(new_n12140));
  inv1 g11947(.a(new_n12138), .O(new_n12141));
  nor2 g11948(.a(new_n12141), .b(new_n12140), .O(new_n12142));
  nor2 g11949(.a(new_n12142), .b(new_n12139), .O(new_n12143));
  nor2 g11950(.a(new_n12143), .b(new_n12130), .O(new_n12144));
  inv1 g11951(.a(new_n12130), .O(new_n12145));
  inv1 g11952(.a(new_n12143), .O(new_n12146));
  nor2 g11953(.a(new_n12146), .b(new_n12145), .O(new_n12147));
  nor2 g11954(.a(new_n12147), .b(new_n12144), .O(new_n12148));
  inv1 g11955(.a(new_n12148), .O(new_n12149));
  nor2 g11956(.a(new_n12149), .b(new_n12117), .O(new_n12150));
  inv1 g11957(.a(new_n12117), .O(new_n12151));
  nor2 g11958(.a(new_n12148), .b(new_n12151), .O(new_n12152));
  nor2 g11959(.a(new_n12152), .b(new_n12150), .O(new_n12153));
  nor2 g11960(.a(new_n12153), .b(new_n12116), .O(new_n12154));
  inv1 g11961(.a(new_n12116), .O(new_n12155));
  inv1 g11962(.a(new_n12153), .O(new_n12156));
  nor2 g11963(.a(new_n12156), .b(new_n12155), .O(new_n12157));
  nor2 g11964(.a(new_n12157), .b(new_n12154), .O(new_n12158));
  inv1 g11965(.a(new_n12158), .O(new_n12159));
  nor2 g11966(.a(new_n12159), .b(new_n12109), .O(new_n12160));
  inv1 g11967(.a(new_n12109), .O(new_n12161));
  nor2 g11968(.a(new_n12158), .b(new_n12161), .O(new_n12162));
  nor2 g11969(.a(new_n12162), .b(new_n12160), .O(new_n12163));
  inv1 g11970(.a(new_n12163), .O(new_n12164));
  nor2 g11971(.a(new_n12164), .b(new_n12108), .O(new_n12165));
  inv1 g11972(.a(new_n12108), .O(new_n12166));
  nor2 g11973(.a(new_n12163), .b(new_n12166), .O(new_n12167));
  nor2 g11974(.a(new_n12167), .b(new_n12165), .O(new_n12168));
  inv1 g11975(.a(new_n12168), .O(new_n12169));
  nor2 g11976(.a(new_n12169), .b(new_n12107), .O(new_n12170));
  inv1 g11977(.a(new_n12107), .O(new_n12171));
  nor2 g11978(.a(new_n12168), .b(new_n12171), .O(new_n12172));
  nor2 g11979(.a(new_n12172), .b(new_n12170), .O(new_n12173));
  inv1 g11980(.a(new_n12173), .O(new_n12174));
  nor2 g11981(.a(new_n12174), .b(new_n12106), .O(new_n12175));
  nor2 g11982(.a(new_n12173), .b(new_n12105), .O(new_n12176));
  nor2 g11983(.a(new_n12176), .b(new_n12175), .O(new_n12177));
  nor2 g11984(.a(new_n11814), .b(new_n11552), .O(new_n12178));
  inv1 g11985(.a(new_n12178), .O(new_n12179));
  nor2 g11986(.a(new_n12179), .b(new_n12177), .O(new_n12180));
  inv1 g11987(.a(new_n12177), .O(new_n12181));
  nor2 g11988(.a(new_n12178), .b(new_n12181), .O(new_n12182));
  nor2 g11989(.a(new_n12182), .b(new_n12180), .O(new_n12183));
  nor2 g11990(.a(new_n11822), .b(new_n11816), .O(new_n12184));
  inv1 g11991(.a(new_n12184), .O(new_n12185));
  nor2 g11992(.a(new_n12185), .b(new_n12183), .O(new_n12186));
  inv1 g11993(.a(new_n12183), .O(new_n12187));
  nor2 g11994(.a(new_n12184), .b(new_n12187), .O(new_n12188));
  nor2 g11995(.a(new_n12188), .b(new_n12186), .O(new_n12189));
  inv1 g11996(.a(new_n12189), .O(\asquared[65] ));
  nor2 g11997(.a(new_n12175), .b(new_n12170), .O(new_n12191));
  nor2 g11998(.a(new_n12103), .b(new_n11923), .O(new_n12192));
  inv1 g11999(.a(new_n12192), .O(new_n12193));
  nor2 g12000(.a(new_n12099), .b(new_n12068), .O(new_n12194));
  nor2 g12001(.a(new_n11920), .b(new_n11857), .O(new_n12195));
  nor2 g12002(.a(new_n12064), .b(new_n12010), .O(new_n12196));
  inv1 g12003(.a(new_n12196), .O(new_n12197));
  nor2 g12004(.a(new_n11914), .b(new_n11864), .O(new_n12198));
  inv1 g12005(.a(new_n12198), .O(new_n12199));
  nor2 g12006(.a(new_n12199), .b(new_n12197), .O(new_n12200));
  nor2 g12007(.a(new_n12198), .b(new_n12196), .O(new_n12201));
  nor2 g12008(.a(new_n12201), .b(new_n12200), .O(new_n12202));
  nor2 g12009(.a(new_n11910), .b(new_n11904), .O(new_n12203));
  nor2 g12010(.a(new_n11902), .b(new_n11896), .O(new_n12204));
  nor2 g12011(.a(new_n12025), .b(new_n12018), .O(new_n12205));
  nor2 g12012(.a(new_n12205), .b(new_n12204), .O(new_n12206));
  inv1 g12013(.a(new_n12204), .O(new_n12207));
  inv1 g12014(.a(new_n12205), .O(new_n12208));
  nor2 g12015(.a(new_n12208), .b(new_n12207), .O(new_n12209));
  nor2 g12016(.a(new_n12209), .b(new_n12206), .O(new_n12210));
  nor2 g12017(.a(new_n12037), .b(new_n12031), .O(new_n12211));
  nor2 g12018(.a(new_n12211), .b(new_n12210), .O(new_n12212));
  inv1 g12019(.a(new_n12210), .O(new_n12213));
  inv1 g12020(.a(new_n12211), .O(new_n12214));
  nor2 g12021(.a(new_n12214), .b(new_n12213), .O(new_n12215));
  nor2 g12022(.a(new_n12215), .b(new_n12212), .O(new_n12216));
  nor2 g12023(.a(new_n11949), .b(new_n11942), .O(new_n12217));
  nor2 g12024(.a(new_n11938), .b(new_n11930), .O(new_n12218));
  nor2 g12025(.a(new_n12218), .b(new_n12217), .O(new_n12219));
  inv1 g12026(.a(new_n12217), .O(new_n12220));
  inv1 g12027(.a(new_n12218), .O(new_n12221));
  nor2 g12028(.a(new_n12221), .b(new_n12220), .O(new_n12222));
  nor2 g12029(.a(new_n12222), .b(new_n12219), .O(new_n12223));
  nor2 g12030(.a(new_n11984), .b(new_n11978), .O(new_n12224));
  nor2 g12031(.a(new_n12224), .b(new_n12223), .O(new_n12225));
  inv1 g12032(.a(new_n12223), .O(new_n12226));
  inv1 g12033(.a(new_n12224), .O(new_n12227));
  nor2 g12034(.a(new_n12227), .b(new_n12226), .O(new_n12228));
  nor2 g12035(.a(new_n12228), .b(new_n12225), .O(new_n12229));
  nor2 g12036(.a(new_n12229), .b(new_n12216), .O(new_n12230));
  inv1 g12037(.a(new_n12216), .O(new_n12231));
  inv1 g12038(.a(new_n12229), .O(new_n12232));
  nor2 g12039(.a(new_n12232), .b(new_n12231), .O(new_n12233));
  nor2 g12040(.a(new_n12233), .b(new_n12230), .O(new_n12234));
  inv1 g12041(.a(new_n12234), .O(new_n12235));
  nor2 g12042(.a(new_n12235), .b(new_n12203), .O(new_n12236));
  inv1 g12043(.a(new_n12203), .O(new_n12237));
  nor2 g12044(.a(new_n12234), .b(new_n12237), .O(new_n12238));
  nor2 g12045(.a(new_n12238), .b(new_n12236), .O(new_n12239));
  nor2 g12046(.a(new_n12239), .b(new_n12202), .O(new_n12240));
  inv1 g12047(.a(new_n12202), .O(new_n12241));
  inv1 g12048(.a(new_n12239), .O(new_n12242));
  nor2 g12049(.a(new_n12242), .b(new_n12241), .O(new_n12243));
  nor2 g12050(.a(new_n12243), .b(new_n12240), .O(new_n12244));
  inv1 g12051(.a(new_n12244), .O(new_n12245));
  nor2 g12052(.a(new_n12245), .b(new_n12195), .O(new_n12246));
  inv1 g12053(.a(new_n12195), .O(new_n12247));
  nor2 g12054(.a(new_n12244), .b(new_n12247), .O(new_n12248));
  nor2 g12055(.a(new_n12248), .b(new_n12246), .O(new_n12249));
  inv1 g12056(.a(new_n12249), .O(new_n12250));
  nor2 g12057(.a(new_n12250), .b(new_n12194), .O(new_n12251));
  inv1 g12058(.a(new_n12194), .O(new_n12252));
  nor2 g12059(.a(new_n12249), .b(new_n12252), .O(new_n12253));
  nor2 g12060(.a(new_n12253), .b(new_n12251), .O(new_n12254));
  nor2 g12061(.a(new_n12254), .b(new_n12193), .O(new_n12255));
  inv1 g12062(.a(new_n12254), .O(new_n12256));
  nor2 g12063(.a(new_n12256), .b(new_n12192), .O(new_n12257));
  nor2 g12064(.a(new_n12257), .b(new_n12255), .O(new_n12258));
  inv1 g12065(.a(new_n12258), .O(new_n12259));
  nor2 g12066(.a(new_n12165), .b(new_n12160), .O(new_n12260));
  nor2 g12067(.a(new_n12052), .b(new_n12044), .O(new_n12261));
  nor2 g12068(.a(new_n11998), .b(new_n11990), .O(new_n12262));
  nor2 g12069(.a(new_n12262), .b(new_n12261), .O(new_n12263));
  inv1 g12070(.a(new_n12261), .O(new_n12264));
  inv1 g12071(.a(new_n12262), .O(new_n12265));
  nor2 g12072(.a(new_n12265), .b(new_n12264), .O(new_n12266));
  nor2 g12073(.a(new_n12266), .b(new_n12263), .O(new_n12267));
  nor2 g12074(.a(new_n11891), .b(new_n11883), .O(new_n12268));
  nor2 g12075(.a(new_n12268), .b(new_n12267), .O(new_n12269));
  inv1 g12076(.a(new_n12267), .O(new_n12270));
  inv1 g12077(.a(new_n12268), .O(new_n12271));
  nor2 g12078(.a(new_n12271), .b(new_n12270), .O(new_n12272));
  nor2 g12079(.a(new_n12272), .b(new_n12269), .O(new_n12273));
  nor2 g12080(.a(new_n12007), .b(new_n12000), .O(new_n12274));
  inv1 g12081(.a(new_n12274), .O(new_n12275));
  nor2 g12082(.a(new_n12275), .b(new_n12273), .O(new_n12276));
  inv1 g12083(.a(new_n12273), .O(new_n12277));
  nor2 g12084(.a(new_n12274), .b(new_n12277), .O(new_n12278));
  nor2 g12085(.a(new_n12278), .b(new_n12276), .O(new_n12279));
  nor2 g12086(.a(new_n12061), .b(new_n12054), .O(new_n12280));
  inv1 g12087(.a(new_n12280), .O(new_n12281));
  nor2 g12088(.a(new_n12281), .b(new_n12279), .O(new_n12282));
  inv1 g12089(.a(new_n12279), .O(new_n12283));
  nor2 g12090(.a(new_n12280), .b(new_n12283), .O(new_n12284));
  nor2 g12091(.a(new_n12284), .b(new_n12282), .O(new_n12285));
  inv1 g12092(.a(new_n12285), .O(new_n12286));
  nor2 g12093(.a(new_n12095), .b(new_n12089), .O(new_n12287));
  nor2 g12094(.a(new_n12287), .b(new_n12286), .O(new_n12288));
  inv1 g12095(.a(new_n12287), .O(new_n12289));
  nor2 g12096(.a(new_n12289), .b(new_n12285), .O(new_n12290));
  nor2 g12097(.a(new_n12290), .b(new_n12288), .O(new_n12291));
  inv1 g12098(.a(new_n12291), .O(new_n12292));
  nor2 g12099(.a(new_n12084), .b(new_n12078), .O(new_n12293));
  inv1 g12100(.a(new_n12293), .O(new_n12294));
  nor2 g12101(.a(new_n11958), .b(new_n11952), .O(new_n12295));
  inv1 g12102(.a(new_n12295), .O(new_n12296));
  nor2 g12103(.a(new_n12296), .b(new_n12294), .O(new_n12297));
  nor2 g12104(.a(new_n12295), .b(new_n12293), .O(new_n12298));
  nor2 g12105(.a(new_n12298), .b(new_n12297), .O(new_n12299));
  inv1 g12106(.a(new_n12299), .O(new_n12300));
  nor2 g12107(.a(new_n11596), .b(new_n196), .O(new_n12301));
  nor2 g12108(.a(new_n12301), .b(new_n11932), .O(new_n12302));
  nor2 g12109(.a(new_n11596), .b(new_n214), .O(new_n12303));
  inv1 g12110(.a(new_n12303), .O(new_n12304));
  nor2 g12111(.a(new_n12304), .b(new_n11720), .O(new_n12305));
  nor2 g12112(.a(new_n12305), .b(new_n12302), .O(new_n12306));
  inv1 g12113(.a(new_n12306), .O(new_n12307));
  nor2 g12114(.a(new_n11974), .b(new_n11967), .O(new_n12308));
  inv1 g12115(.a(new_n12308), .O(new_n12309));
  nor2 g12116(.a(new_n12309), .b(new_n12307), .O(new_n12310));
  nor2 g12117(.a(new_n12308), .b(new_n12306), .O(new_n12311));
  nor2 g12118(.a(new_n12311), .b(new_n12310), .O(new_n12312));
  inv1 g12119(.a(new_n12312), .O(new_n12313));
  nor2 g12120(.a(new_n7294), .b(new_n800), .O(new_n12314));
  nor2 g12121(.a(new_n7537), .b(new_n699), .O(new_n12315));
  nor2 g12122(.a(new_n12315), .b(new_n12314), .O(new_n12316));
  nor2 g12123(.a(new_n11964), .b(new_n10862), .O(new_n12317));
  nor2 g12124(.a(new_n12317), .b(new_n12316), .O(new_n12318));
  nor2 g12125(.a(new_n12318), .b(new_n9597), .O(new_n12319));
  inv1 g12126(.a(new_n12318), .O(new_n12320));
  nor2 g12127(.a(new_n12320), .b(new_n9596), .O(new_n12321));
  nor2 g12128(.a(new_n12321), .b(new_n12319), .O(new_n12322));
  nor2 g12129(.a(new_n8026), .b(new_n613), .O(new_n12323));
  nor2 g12130(.a(new_n6570), .b(new_n1086), .O(new_n12324));
  nor2 g12131(.a(new_n12324), .b(new_n12323), .O(new_n12325));
  inv1 g12132(.a(new_n12323), .O(new_n12326));
  inv1 g12133(.a(new_n12324), .O(new_n12327));
  nor2 g12134(.a(new_n12327), .b(new_n12326), .O(new_n12328));
  nor2 g12135(.a(new_n12328), .b(new_n12325), .O(new_n12329));
  nor2 g12136(.a(new_n12329), .b(new_n11886), .O(new_n12330));
  inv1 g12137(.a(new_n12329), .O(new_n12331));
  nor2 g12138(.a(new_n12331), .b(new_n11885), .O(new_n12332));
  nor2 g12139(.a(new_n12332), .b(new_n12330), .O(new_n12333));
  nor2 g12140(.a(new_n12333), .b(new_n12322), .O(new_n12334));
  inv1 g12141(.a(new_n12322), .O(new_n12335));
  inv1 g12142(.a(new_n12333), .O(new_n12336));
  nor2 g12143(.a(new_n12336), .b(new_n12335), .O(new_n12337));
  nor2 g12144(.a(new_n12337), .b(new_n12334), .O(new_n12338));
  inv1 g12145(.a(new_n12338), .O(new_n12339));
  nor2 g12146(.a(new_n12339), .b(new_n12313), .O(new_n12340));
  nor2 g12147(.a(new_n12338), .b(new_n12312), .O(new_n12341));
  nor2 g12148(.a(new_n12341), .b(new_n12340), .O(new_n12342));
  inv1 g12149(.a(new_n12342), .O(new_n12343));
  nor2 g12150(.a(new_n12343), .b(new_n12300), .O(new_n12344));
  nor2 g12151(.a(new_n12342), .b(new_n12299), .O(new_n12345));
  nor2 g12152(.a(new_n12345), .b(new_n12344), .O(new_n12346));
  inv1 g12153(.a(new_n12346), .O(new_n12347));
  nor2 g12154(.a(new_n12347), .b(new_n12292), .O(new_n12348));
  nor2 g12155(.a(new_n12346), .b(new_n12291), .O(new_n12349));
  nor2 g12156(.a(new_n12349), .b(new_n12348), .O(new_n12350));
  inv1 g12157(.a(new_n12350), .O(new_n12351));
  nor2 g12158(.a(new_n12351), .b(new_n12260), .O(new_n12352));
  inv1 g12159(.a(new_n12260), .O(new_n12353));
  nor2 g12160(.a(new_n12350), .b(new_n12353), .O(new_n12354));
  nor2 g12161(.a(new_n12354), .b(new_n12352), .O(new_n12355));
  inv1 g12162(.a(new_n12355), .O(new_n12356));
  nor2 g12163(.a(new_n11839), .b(new_n11833), .O(new_n12357));
  inv1 g12164(.a(new_n12357), .O(new_n12358));
  nor2 g12165(.a(new_n12129), .b(new_n12123), .O(new_n12359));
  inv1 g12166(.a(new_n12359), .O(new_n12360));
  nor2 g12167(.a(new_n12360), .b(new_n12358), .O(new_n12361));
  nor2 g12168(.a(new_n12359), .b(new_n12357), .O(new_n12362));
  nor2 g12169(.a(new_n12362), .b(new_n12361), .O(new_n12363));
  nor2 g12170(.a(new_n12142), .b(new_n12136), .O(new_n12364));
  inv1 g12171(.a(new_n12364), .O(new_n12365));
  nor2 g12172(.a(new_n12365), .b(new_n12363), .O(new_n12366));
  inv1 g12173(.a(new_n12363), .O(new_n12367));
  nor2 g12174(.a(new_n12364), .b(new_n12367), .O(new_n12368));
  nor2 g12175(.a(new_n12368), .b(new_n12366), .O(new_n12369));
  inv1 g12176(.a(new_n12369), .O(new_n12370));
  nor2 g12177(.a(new_n12150), .b(new_n12147), .O(new_n12371));
  nor2 g12178(.a(new_n11851), .b(new_n11845), .O(new_n12372));
  nor2 g12179(.a(new_n12372), .b(new_n12371), .O(new_n12373));
  inv1 g12180(.a(new_n12371), .O(new_n12374));
  inv1 g12181(.a(new_n12372), .O(new_n12375));
  nor2 g12182(.a(new_n12375), .b(new_n12374), .O(new_n12376));
  nor2 g12183(.a(new_n12376), .b(new_n12373), .O(new_n12377));
  inv1 g12184(.a(new_n12377), .O(new_n12378));
  nor2 g12185(.a(new_n12378), .b(new_n12370), .O(new_n12379));
  nor2 g12186(.a(new_n12377), .b(new_n12369), .O(new_n12380));
  nor2 g12187(.a(new_n12380), .b(new_n12379), .O(new_n12381));
  inv1 g12188(.a(new_n12381), .O(new_n12382));
  nor2 g12189(.a(new_n12157), .b(new_n12115), .O(new_n12383));
  nor2 g12190(.a(new_n10468), .b(new_n229), .O(new_n12384));
  inv1 g12191(.a(new_n12384), .O(new_n12385));
  nor2 g12192(.a(new_n10320), .b(new_n257), .O(new_n12386));
  nor2 g12193(.a(new_n9873), .b(new_n295), .O(new_n12387));
  nor2 g12194(.a(new_n12387), .b(new_n12386), .O(new_n12388));
  nor2 g12195(.a(new_n10320), .b(new_n295), .O(new_n12389));
  inv1 g12196(.a(new_n12389), .O(new_n12390));
  nor2 g12197(.a(new_n12390), .b(new_n12038), .O(new_n12391));
  nor2 g12198(.a(new_n12391), .b(new_n12388), .O(new_n12392));
  nor2 g12199(.a(new_n12392), .b(new_n12385), .O(new_n12393));
  inv1 g12200(.a(new_n12392), .O(new_n12394));
  nor2 g12201(.a(new_n12394), .b(new_n12384), .O(new_n12395));
  nor2 g12202(.a(new_n12395), .b(new_n12393), .O(new_n12396));
  nor2 g12203(.a(new_n9658), .b(new_n322), .O(new_n12397));
  inv1 g12204(.a(new_n12397), .O(new_n12398));
  nor2 g12205(.a(new_n5796), .b(new_n1425), .O(new_n12399));
  nor2 g12206(.a(new_n12399), .b(new_n12046), .O(new_n12400));
  inv1 g12207(.a(new_n12043), .O(new_n12401));
  nor2 g12208(.a(new_n5796), .b(new_n1493), .O(new_n12402));
  inv1 g12209(.a(new_n12402), .O(new_n12403));
  nor2 g12210(.a(new_n12403), .b(new_n12401), .O(new_n12404));
  nor2 g12211(.a(new_n12404), .b(new_n12400), .O(new_n12405));
  nor2 g12212(.a(new_n12405), .b(new_n12398), .O(new_n12406));
  inv1 g12213(.a(new_n12405), .O(new_n12407));
  nor2 g12214(.a(new_n12407), .b(new_n12397), .O(new_n12408));
  nor2 g12215(.a(new_n12408), .b(new_n12406), .O(new_n12409));
  nor2 g12216(.a(new_n11877), .b(new_n11870), .O(new_n12410));
  nor2 g12217(.a(new_n12410), .b(new_n12409), .O(new_n12411));
  inv1 g12218(.a(new_n12409), .O(new_n12412));
  inv1 g12219(.a(new_n12410), .O(new_n12413));
  nor2 g12220(.a(new_n12413), .b(new_n12412), .O(new_n12414));
  nor2 g12221(.a(new_n12414), .b(new_n12411), .O(new_n12415));
  inv1 g12222(.a(new_n12415), .O(new_n12416));
  nor2 g12223(.a(new_n12416), .b(new_n12396), .O(new_n12417));
  inv1 g12224(.a(new_n12396), .O(new_n12418));
  nor2 g12225(.a(new_n12415), .b(new_n12418), .O(new_n12419));
  nor2 g12226(.a(new_n12419), .b(new_n12417), .O(new_n12420));
  inv1 g12227(.a(new_n12420), .O(new_n12421));
  nor2 g12228(.a(new_n8476), .b(new_n502), .O(new_n12422));
  nor2 g12229(.a(new_n12422), .b(new_n11943), .O(new_n12423));
  inv1 g12230(.a(new_n12422), .O(new_n12424));
  nor2 g12231(.a(new_n12424), .b(new_n11944), .O(new_n12425));
  nor2 g12232(.a(new_n12425), .b(new_n12423), .O(new_n12426));
  inv1 g12233(.a(new_n12426), .O(new_n12427));
  nor2 g12234(.a(new_n12427), .b(new_n11993), .O(new_n12428));
  nor2 g12235(.a(new_n12426), .b(new_n11992), .O(new_n12429));
  nor2 g12236(.a(new_n12429), .b(new_n12428), .O(new_n12430));
  inv1 g12237(.a(new_n12430), .O(new_n12431));
  nor2 g12238(.a(new_n3722), .b(new_n2660), .O(new_n12432));
  inv1 g12239(.a(new_n12432), .O(new_n12433));
  nor2 g12240(.a(new_n3231), .b(new_n3057), .O(new_n12434));
  nor2 g12241(.a(new_n12434), .b(new_n11968), .O(new_n12435));
  inv1 g12242(.a(new_n11965), .O(new_n12436));
  nor2 g12243(.a(new_n3533), .b(new_n3057), .O(new_n12437));
  inv1 g12244(.a(new_n12437), .O(new_n12438));
  nor2 g12245(.a(new_n12438), .b(new_n12436), .O(new_n12439));
  nor2 g12246(.a(new_n12439), .b(new_n12435), .O(new_n12440));
  nor2 g12247(.a(new_n12440), .b(new_n12433), .O(new_n12441));
  inv1 g12248(.a(new_n12440), .O(new_n12442));
  nor2 g12249(.a(new_n12442), .b(new_n12432), .O(new_n12443));
  nor2 g12250(.a(new_n12443), .b(new_n12441), .O(new_n12444));
  nor2 g12251(.a(new_n12444), .b(new_n12431), .O(new_n12445));
  inv1 g12252(.a(new_n12444), .O(new_n12446));
  nor2 g12253(.a(new_n12446), .b(new_n12430), .O(new_n12447));
  nor2 g12254(.a(new_n12447), .b(new_n12445), .O(new_n12448));
  inv1 g12255(.a(new_n12448), .O(new_n12449));
  nor2 g12256(.a(new_n6893), .b(new_n941), .O(new_n12450));
  inv1 g12257(.a(new_n12450), .O(new_n12451));
  nor2 g12258(.a(new_n11186), .b(new_n203), .O(new_n12452));
  inv1 g12259(.a(new_n12452), .O(new_n12453));
  nor2 g12260(.a(new_n12453), .b(new_n3231), .O(new_n12454));
  nor2 g12261(.a(new_n12452), .b(\a[33] ), .O(new_n12455));
  nor2 g12262(.a(new_n12455), .b(new_n12454), .O(new_n12456));
  nor2 g12263(.a(new_n12456), .b(new_n12451), .O(new_n12457));
  inv1 g12264(.a(new_n12456), .O(new_n12458));
  nor2 g12265(.a(new_n12458), .b(new_n12450), .O(new_n12459));
  nor2 g12266(.a(new_n12459), .b(new_n12457), .O(new_n12460));
  nor2 g12267(.a(new_n12460), .b(new_n12449), .O(new_n12461));
  inv1 g12268(.a(new_n12460), .O(new_n12462));
  nor2 g12269(.a(new_n12462), .b(new_n12448), .O(new_n12463));
  nor2 g12270(.a(new_n12463), .b(new_n12461), .O(new_n12464));
  inv1 g12271(.a(new_n12464), .O(new_n12465));
  nor2 g12272(.a(new_n12465), .b(new_n12421), .O(new_n12466));
  nor2 g12273(.a(new_n12464), .b(new_n12420), .O(new_n12467));
  nor2 g12274(.a(new_n12467), .b(new_n12466), .O(new_n12468));
  inv1 g12275(.a(new_n12468), .O(new_n12469));
  nor2 g12276(.a(new_n4425), .b(new_n2121), .O(new_n12470));
  inv1 g12277(.a(new_n12470), .O(new_n12471));
  nor2 g12278(.a(new_n4093), .b(new_n2433), .O(new_n12472));
  nor2 g12279(.a(new_n4366), .b(new_n2184), .O(new_n12473));
  nor2 g12280(.a(new_n12473), .b(new_n12472), .O(new_n12474));
  nor2 g12281(.a(new_n4366), .b(new_n2433), .O(new_n12475));
  inv1 g12282(.a(new_n12475), .O(new_n12476));
  nor2 g12283(.a(new_n12476), .b(new_n11988), .O(new_n12477));
  nor2 g12284(.a(new_n12477), .b(new_n12474), .O(new_n12478));
  nor2 g12285(.a(new_n12478), .b(new_n12471), .O(new_n12479));
  inv1 g12286(.a(new_n12478), .O(new_n12480));
  nor2 g12287(.a(new_n12480), .b(new_n12470), .O(new_n12481));
  nor2 g12288(.a(new_n12481), .b(new_n12479), .O(new_n12482));
  inv1 g12289(.a(new_n12482), .O(new_n12483));
  nor2 g12290(.a(new_n5178), .b(new_n1647), .O(new_n12484));
  inv1 g12291(.a(new_n12484), .O(new_n12485));
  nor2 g12292(.a(new_n4954), .b(new_n1736), .O(new_n12486));
  nor2 g12293(.a(new_n12486), .b(new_n12019), .O(new_n12487));
  inv1 g12294(.a(new_n12016), .O(new_n12488));
  nor2 g12295(.a(new_n4954), .b(new_n1903), .O(new_n12489));
  inv1 g12296(.a(new_n12489), .O(new_n12490));
  nor2 g12297(.a(new_n12490), .b(new_n12488), .O(new_n12491));
  nor2 g12298(.a(new_n12491), .b(new_n12487), .O(new_n12492));
  nor2 g12299(.a(new_n12492), .b(new_n12485), .O(new_n12493));
  inv1 g12300(.a(new_n12492), .O(new_n12494));
  nor2 g12301(.a(new_n12494), .b(new_n12484), .O(new_n12495));
  nor2 g12302(.a(new_n12495), .b(new_n12493), .O(new_n12496));
  nor2 g12303(.a(new_n9156), .b(new_n363), .O(new_n12497));
  inv1 g12304(.a(new_n12497), .O(new_n12498));
  nor2 g12305(.a(new_n8946), .b(new_n438), .O(new_n12499));
  nor2 g12306(.a(new_n5971), .b(new_n1297), .O(new_n12500));
  nor2 g12307(.a(new_n12500), .b(new_n12499), .O(new_n12501));
  inv1 g12308(.a(new_n12499), .O(new_n12502));
  inv1 g12309(.a(new_n12500), .O(new_n12503));
  nor2 g12310(.a(new_n12503), .b(new_n12502), .O(new_n12504));
  nor2 g12311(.a(new_n12504), .b(new_n12501), .O(new_n12505));
  nor2 g12312(.a(new_n12505), .b(new_n12498), .O(new_n12506));
  inv1 g12313(.a(new_n12505), .O(new_n12507));
  nor2 g12314(.a(new_n12507), .b(new_n12497), .O(new_n12508));
  nor2 g12315(.a(new_n12508), .b(new_n12506), .O(new_n12509));
  nor2 g12316(.a(new_n12509), .b(new_n12496), .O(new_n12510));
  inv1 g12317(.a(new_n12496), .O(new_n12511));
  inv1 g12318(.a(new_n12509), .O(new_n12512));
  nor2 g12319(.a(new_n12512), .b(new_n12511), .O(new_n12513));
  nor2 g12320(.a(new_n12513), .b(new_n12510), .O(new_n12514));
  nor2 g12321(.a(new_n12514), .b(new_n12483), .O(new_n12515));
  inv1 g12322(.a(new_n12514), .O(new_n12516));
  nor2 g12323(.a(new_n12516), .b(new_n12482), .O(new_n12517));
  nor2 g12324(.a(new_n12517), .b(new_n12515), .O(new_n12518));
  inv1 g12325(.a(new_n12518), .O(new_n12519));
  nor2 g12326(.a(new_n12519), .b(new_n12469), .O(new_n12520));
  nor2 g12327(.a(new_n12518), .b(new_n12468), .O(new_n12521));
  nor2 g12328(.a(new_n12521), .b(new_n12520), .O(new_n12522));
  inv1 g12329(.a(new_n12522), .O(new_n12523));
  nor2 g12330(.a(new_n12523), .b(new_n12383), .O(new_n12524));
  inv1 g12331(.a(new_n12383), .O(new_n12525));
  nor2 g12332(.a(new_n12522), .b(new_n12525), .O(new_n12526));
  nor2 g12333(.a(new_n12526), .b(new_n12524), .O(new_n12527));
  inv1 g12334(.a(new_n12527), .O(new_n12528));
  nor2 g12335(.a(new_n12528), .b(new_n12382), .O(new_n12529));
  nor2 g12336(.a(new_n12527), .b(new_n12381), .O(new_n12530));
  nor2 g12337(.a(new_n12530), .b(new_n12529), .O(new_n12531));
  inv1 g12338(.a(new_n12531), .O(new_n12532));
  nor2 g12339(.a(new_n12532), .b(new_n12356), .O(new_n12533));
  nor2 g12340(.a(new_n12531), .b(new_n12355), .O(new_n12534));
  nor2 g12341(.a(new_n12534), .b(new_n12533), .O(new_n12535));
  inv1 g12342(.a(new_n12535), .O(new_n12536));
  nor2 g12343(.a(new_n12536), .b(new_n12259), .O(new_n12537));
  nor2 g12344(.a(new_n12535), .b(new_n12258), .O(new_n12538));
  nor2 g12345(.a(new_n12538), .b(new_n12537), .O(new_n12539));
  inv1 g12346(.a(new_n12539), .O(new_n12540));
  nor2 g12347(.a(new_n12540), .b(new_n12191), .O(new_n12541));
  inv1 g12348(.a(new_n12191), .O(new_n12542));
  nor2 g12349(.a(new_n12539), .b(new_n12542), .O(new_n12543));
  nor2 g12350(.a(new_n12543), .b(new_n12541), .O(new_n12544));
  inv1 g12351(.a(new_n12544), .O(new_n12545));
  nor2 g12352(.a(new_n12188), .b(new_n12180), .O(new_n12546));
  nor2 g12353(.a(new_n12546), .b(new_n12545), .O(new_n12547));
  inv1 g12354(.a(new_n12546), .O(new_n12548));
  nor2 g12355(.a(new_n12548), .b(new_n12544), .O(new_n12549));
  nor2 g12356(.a(new_n12549), .b(new_n12547), .O(new_n12550));
  inv1 g12357(.a(new_n12550), .O(\asquared[66] ));
  nor2 g12358(.a(new_n12537), .b(new_n12257), .O(new_n12552));
  nor2 g12359(.a(new_n12251), .b(new_n12246), .O(new_n12553));
  inv1 g12360(.a(new_n12553), .O(new_n12554));
  nor2 g12361(.a(new_n12529), .b(new_n12524), .O(new_n12555));
  inv1 g12362(.a(new_n12555), .O(new_n12556));
  nor2 g12363(.a(new_n12556), .b(new_n12554), .O(new_n12557));
  nor2 g12364(.a(new_n12555), .b(new_n12553), .O(new_n12558));
  nor2 g12365(.a(new_n12558), .b(new_n12557), .O(new_n12559));
  inv1 g12366(.a(new_n12559), .O(new_n12560));
  nor2 g12367(.a(new_n12243), .b(new_n12201), .O(new_n12561));
  nor2 g12368(.a(new_n9156), .b(new_n438), .O(new_n12562));
  inv1 g12369(.a(new_n12562), .O(new_n12563));
  nor2 g12370(.a(new_n4682), .b(new_n2121), .O(new_n12564));
  nor2 g12371(.a(new_n12564), .b(new_n12489), .O(new_n12565));
  nor2 g12372(.a(new_n4954), .b(new_n2121), .O(new_n12566));
  inv1 g12373(.a(new_n12566), .O(new_n12567));
  nor2 g12374(.a(new_n12567), .b(new_n12020), .O(new_n12568));
  nor2 g12375(.a(new_n12568), .b(new_n12565), .O(new_n12569));
  nor2 g12376(.a(new_n12569), .b(new_n12563), .O(new_n12570));
  inv1 g12377(.a(new_n12569), .O(new_n12571));
  nor2 g12378(.a(new_n12571), .b(new_n12562), .O(new_n12572));
  nor2 g12379(.a(new_n12572), .b(new_n12570), .O(new_n12573));
  inv1 g12380(.a(new_n12573), .O(new_n12574));
  nor2 g12381(.a(new_n5393), .b(new_n1647), .O(new_n12575));
  nor2 g12382(.a(new_n9658), .b(new_n363), .O(new_n12576));
  nor2 g12383(.a(new_n5178), .b(new_n1736), .O(new_n12577));
  nor2 g12384(.a(new_n12577), .b(new_n12576), .O(new_n12578));
  nor2 g12385(.a(new_n9658), .b(new_n1736), .O(new_n12579));
  inv1 g12386(.a(new_n12579), .O(new_n12580));
  nor2 g12387(.a(new_n12580), .b(new_n7637), .O(new_n12581));
  nor2 g12388(.a(new_n12581), .b(new_n12578), .O(new_n12582));
  inv1 g12389(.a(new_n12582), .O(new_n12583));
  nor2 g12390(.a(new_n12583), .b(new_n12575), .O(new_n12584));
  inv1 g12391(.a(new_n12575), .O(new_n12585));
  nor2 g12392(.a(new_n12582), .b(new_n12585), .O(new_n12586));
  nor2 g12393(.a(new_n12586), .b(new_n12584), .O(new_n12587));
  nor2 g12394(.a(new_n6274), .b(new_n1297), .O(new_n12588));
  inv1 g12395(.a(new_n12588), .O(new_n12589));
  nor2 g12396(.a(new_n5971), .b(new_n1425), .O(new_n12590));
  nor2 g12397(.a(new_n12590), .b(new_n12402), .O(new_n12591));
  inv1 g12398(.a(new_n12399), .O(new_n12592));
  nor2 g12399(.a(new_n5971), .b(new_n1493), .O(new_n12593));
  inv1 g12400(.a(new_n12593), .O(new_n12594));
  nor2 g12401(.a(new_n12594), .b(new_n12592), .O(new_n12595));
  nor2 g12402(.a(new_n12595), .b(new_n12591), .O(new_n12596));
  nor2 g12403(.a(new_n12596), .b(new_n12589), .O(new_n12597));
  inv1 g12404(.a(new_n12596), .O(new_n12598));
  nor2 g12405(.a(new_n12598), .b(new_n12588), .O(new_n12599));
  nor2 g12406(.a(new_n12599), .b(new_n12597), .O(new_n12600));
  nor2 g12407(.a(new_n12600), .b(new_n12587), .O(new_n12601));
  inv1 g12408(.a(new_n12587), .O(new_n12602));
  inv1 g12409(.a(new_n12600), .O(new_n12603));
  nor2 g12410(.a(new_n12603), .b(new_n12602), .O(new_n12604));
  nor2 g12411(.a(new_n12604), .b(new_n12601), .O(new_n12605));
  nor2 g12412(.a(new_n12605), .b(new_n12574), .O(new_n12606));
  inv1 g12413(.a(new_n12605), .O(new_n12607));
  nor2 g12414(.a(new_n12607), .b(new_n12573), .O(new_n12608));
  nor2 g12415(.a(new_n12608), .b(new_n12606), .O(new_n12609));
  inv1 g12416(.a(new_n12609), .O(new_n12610));
  nor2 g12417(.a(new_n7294), .b(new_n847), .O(new_n12611));
  nor2 g12418(.a(new_n12611), .b(new_n8986), .O(new_n12612));
  nor2 g12419(.a(new_n7294), .b(new_n941), .O(new_n12613));
  inv1 g12420(.a(new_n12613), .O(new_n12614));
  nor2 g12421(.a(new_n12614), .b(new_n9597), .O(new_n12615));
  nor2 g12422(.a(new_n12615), .b(new_n12612), .O(new_n12616));
  nor2 g12423(.a(new_n12616), .b(new_n12438), .O(new_n12617));
  inv1 g12424(.a(new_n12616), .O(new_n12618));
  nor2 g12425(.a(new_n12618), .b(new_n12437), .O(new_n12619));
  nor2 g12426(.a(new_n12619), .b(new_n12617), .O(new_n12620));
  inv1 g12427(.a(new_n12620), .O(new_n12621));
  nor2 g12428(.a(new_n6893), .b(new_n1086), .O(new_n12622));
  nor2 g12429(.a(new_n8170), .b(new_n613), .O(new_n12623));
  nor2 g12430(.a(new_n12623), .b(new_n10861), .O(new_n12624));
  nor2 g12431(.a(new_n8170), .b(new_n800), .O(new_n12625));
  inv1 g12432(.a(new_n12625), .O(new_n12626));
  nor2 g12433(.a(new_n12626), .b(new_n11696), .O(new_n12627));
  nor2 g12434(.a(new_n12627), .b(new_n12624), .O(new_n12628));
  inv1 g12435(.a(new_n12628), .O(new_n12629));
  nor2 g12436(.a(new_n12629), .b(new_n12622), .O(new_n12630));
  inv1 g12437(.a(new_n12622), .O(new_n12631));
  nor2 g12438(.a(new_n12628), .b(new_n12631), .O(new_n12632));
  nor2 g12439(.a(new_n12632), .b(new_n12630), .O(new_n12633));
  nor2 g12440(.a(new_n8026), .b(new_n699), .O(new_n12634));
  inv1 g12441(.a(new_n12634), .O(new_n12635));
  nor2 g12442(.a(new_n3722), .b(new_n2826), .O(new_n12636));
  nor2 g12443(.a(new_n3870), .b(new_n2660), .O(new_n12637));
  nor2 g12444(.a(new_n12637), .b(new_n12636), .O(new_n12638));
  nor2 g12445(.a(new_n3870), .b(new_n2826), .O(new_n12639));
  inv1 g12446(.a(new_n12639), .O(new_n12640));
  nor2 g12447(.a(new_n12640), .b(new_n12433), .O(new_n12641));
  nor2 g12448(.a(new_n12641), .b(new_n12638), .O(new_n12642));
  nor2 g12449(.a(new_n12642), .b(new_n12635), .O(new_n12643));
  inv1 g12450(.a(new_n12642), .O(new_n12644));
  nor2 g12451(.a(new_n12644), .b(new_n12634), .O(new_n12645));
  nor2 g12452(.a(new_n12645), .b(new_n12643), .O(new_n12646));
  nor2 g12453(.a(new_n12646), .b(new_n12633), .O(new_n12647));
  inv1 g12454(.a(new_n12633), .O(new_n12648));
  inv1 g12455(.a(new_n12646), .O(new_n12649));
  nor2 g12456(.a(new_n12649), .b(new_n12648), .O(new_n12650));
  nor2 g12457(.a(new_n12650), .b(new_n12647), .O(new_n12651));
  nor2 g12458(.a(new_n12651), .b(new_n12621), .O(new_n12652));
  inv1 g12459(.a(new_n12651), .O(new_n12653));
  nor2 g12460(.a(new_n12653), .b(new_n12620), .O(new_n12654));
  nor2 g12461(.a(new_n12654), .b(new_n12652), .O(new_n12655));
  inv1 g12462(.a(new_n12655), .O(new_n12656));
  nor2 g12463(.a(new_n12656), .b(new_n12610), .O(new_n12657));
  nor2 g12464(.a(new_n12655), .b(new_n12609), .O(new_n12658));
  nor2 g12465(.a(new_n12658), .b(new_n12657), .O(new_n12659));
  inv1 g12466(.a(new_n12659), .O(new_n12660));
  nor2 g12467(.a(new_n8946), .b(new_n502), .O(new_n12661));
  inv1 g12468(.a(new_n12661), .O(new_n12662));
  nor2 g12469(.a(new_n6570), .b(new_n1199), .O(new_n12663));
  nor2 g12470(.a(new_n8476), .b(new_n569), .O(new_n12664));
  nor2 g12471(.a(new_n12664), .b(new_n12663), .O(new_n12665));
  inv1 g12472(.a(new_n12663), .O(new_n12666));
  inv1 g12473(.a(new_n12664), .O(new_n12667));
  nor2 g12474(.a(new_n12667), .b(new_n12666), .O(new_n12668));
  nor2 g12475(.a(new_n12668), .b(new_n12665), .O(new_n12669));
  nor2 g12476(.a(new_n12669), .b(new_n12662), .O(new_n12670));
  inv1 g12477(.a(new_n12669), .O(new_n12671));
  nor2 g12478(.a(new_n12671), .b(new_n12661), .O(new_n12672));
  nor2 g12479(.a(new_n12672), .b(new_n12670), .O(new_n12673));
  inv1 g12480(.a(new_n12673), .O(new_n12674));
  nor2 g12481(.a(new_n11596), .b(new_n203), .O(new_n12675));
  nor2 g12482(.a(new_n10895), .b(new_n229), .O(new_n12676));
  nor2 g12483(.a(new_n11186), .b(new_n214), .O(new_n12677));
  nor2 g12484(.a(new_n12677), .b(new_n12676), .O(new_n12678));
  nor2 g12485(.a(new_n11186), .b(new_n229), .O(new_n12679));
  inv1 g12486(.a(new_n12679), .O(new_n12680));
  nor2 g12487(.a(new_n12680), .b(new_n11933), .O(new_n12681));
  nor2 g12488(.a(new_n12681), .b(new_n12678), .O(new_n12682));
  inv1 g12489(.a(new_n12682), .O(new_n12683));
  nor2 g12490(.a(new_n12683), .b(new_n12675), .O(new_n12684));
  inv1 g12491(.a(new_n12675), .O(new_n12685));
  nor2 g12492(.a(new_n12682), .b(new_n12685), .O(new_n12686));
  nor2 g12493(.a(new_n12686), .b(new_n12684), .O(new_n12687));
  nor2 g12494(.a(new_n4425), .b(new_n2184), .O(new_n12688));
  inv1 g12495(.a(new_n12688), .O(new_n12689));
  nor2 g12496(.a(new_n4093), .b(new_n2506), .O(new_n12690));
  nor2 g12497(.a(new_n12690), .b(new_n12475), .O(new_n12691));
  inv1 g12498(.a(new_n12472), .O(new_n12692));
  nor2 g12499(.a(new_n4366), .b(new_n2506), .O(new_n12693));
  inv1 g12500(.a(new_n12693), .O(new_n12694));
  nor2 g12501(.a(new_n12694), .b(new_n12692), .O(new_n12695));
  nor2 g12502(.a(new_n12695), .b(new_n12691), .O(new_n12696));
  nor2 g12503(.a(new_n12696), .b(new_n12689), .O(new_n12697));
  inv1 g12504(.a(new_n12696), .O(new_n12698));
  nor2 g12505(.a(new_n12698), .b(new_n12688), .O(new_n12699));
  nor2 g12506(.a(new_n12699), .b(new_n12697), .O(new_n12700));
  nor2 g12507(.a(new_n12700), .b(new_n12687), .O(new_n12701));
  inv1 g12508(.a(new_n12687), .O(new_n12702));
  inv1 g12509(.a(new_n12700), .O(new_n12703));
  nor2 g12510(.a(new_n12703), .b(new_n12702), .O(new_n12704));
  nor2 g12511(.a(new_n12704), .b(new_n12701), .O(new_n12705));
  nor2 g12512(.a(new_n12705), .b(new_n12674), .O(new_n12706));
  inv1 g12513(.a(new_n12705), .O(new_n12707));
  nor2 g12514(.a(new_n12707), .b(new_n12673), .O(new_n12708));
  nor2 g12515(.a(new_n12708), .b(new_n12706), .O(new_n12709));
  inv1 g12516(.a(new_n12709), .O(new_n12710));
  nor2 g12517(.a(new_n12710), .b(new_n12660), .O(new_n12711));
  nor2 g12518(.a(new_n12709), .b(new_n12659), .O(new_n12712));
  nor2 g12519(.a(new_n12712), .b(new_n12711), .O(new_n12713));
  inv1 g12520(.a(new_n12713), .O(new_n12714));
  nor2 g12521(.a(new_n12714), .b(new_n12561), .O(new_n12715));
  inv1 g12522(.a(new_n12561), .O(new_n12716));
  nor2 g12523(.a(new_n12713), .b(new_n12716), .O(new_n12717));
  nor2 g12524(.a(new_n12717), .b(new_n12715), .O(new_n12718));
  inv1 g12525(.a(new_n12718), .O(new_n12719));
  nor2 g12526(.a(new_n12215), .b(new_n12209), .O(new_n12720));
  inv1 g12527(.a(new_n12720), .O(new_n12721));
  nor2 g12528(.a(new_n12228), .b(new_n12222), .O(new_n12722));
  inv1 g12529(.a(new_n12722), .O(new_n12723));
  nor2 g12530(.a(new_n12723), .b(new_n12721), .O(new_n12724));
  nor2 g12531(.a(new_n12722), .b(new_n12720), .O(new_n12725));
  nor2 g12532(.a(new_n12725), .b(new_n12724), .O(new_n12726));
  nor2 g12533(.a(new_n12272), .b(new_n12266), .O(new_n12727));
  inv1 g12534(.a(new_n12727), .O(new_n12728));
  nor2 g12535(.a(new_n12728), .b(new_n12726), .O(new_n12729));
  inv1 g12536(.a(new_n12726), .O(new_n12730));
  nor2 g12537(.a(new_n12727), .b(new_n12730), .O(new_n12731));
  nor2 g12538(.a(new_n12731), .b(new_n12729), .O(new_n12732));
  inv1 g12539(.a(new_n12732), .O(new_n12733));
  nor2 g12540(.a(new_n12236), .b(new_n12233), .O(new_n12734));
  nor2 g12541(.a(new_n12284), .b(new_n12278), .O(new_n12735));
  nor2 g12542(.a(new_n12735), .b(new_n12734), .O(new_n12736));
  inv1 g12543(.a(new_n12734), .O(new_n12737));
  inv1 g12544(.a(new_n12735), .O(new_n12738));
  nor2 g12545(.a(new_n12738), .b(new_n12737), .O(new_n12739));
  nor2 g12546(.a(new_n12739), .b(new_n12736), .O(new_n12740));
  inv1 g12547(.a(new_n12740), .O(new_n12741));
  nor2 g12548(.a(new_n12741), .b(new_n12733), .O(new_n12742));
  nor2 g12549(.a(new_n12740), .b(new_n12732), .O(new_n12743));
  nor2 g12550(.a(new_n12743), .b(new_n12742), .O(new_n12744));
  inv1 g12551(.a(new_n12744), .O(new_n12745));
  nor2 g12552(.a(new_n12745), .b(new_n12719), .O(new_n12746));
  nor2 g12553(.a(new_n12744), .b(new_n12718), .O(new_n12747));
  nor2 g12554(.a(new_n12747), .b(new_n12746), .O(new_n12748));
  inv1 g12555(.a(new_n12748), .O(new_n12749));
  nor2 g12556(.a(new_n12749), .b(new_n12560), .O(new_n12750));
  nor2 g12557(.a(new_n12748), .b(new_n12559), .O(new_n12751));
  nor2 g12558(.a(new_n12751), .b(new_n12750), .O(new_n12752));
  inv1 g12559(.a(new_n12752), .O(new_n12753));
  nor2 g12560(.a(new_n12533), .b(new_n12352), .O(new_n12754));
  nor2 g12561(.a(new_n12379), .b(new_n12373), .O(new_n12755));
  nor2 g12562(.a(new_n12368), .b(new_n12362), .O(new_n12756));
  inv1 g12563(.a(new_n12756), .O(new_n12757));
  nor2 g12564(.a(new_n12340), .b(new_n12334), .O(new_n12758));
  nor2 g12565(.a(new_n12310), .b(new_n12305), .O(new_n12759));
  inv1 g12566(.a(new_n12759), .O(new_n12760));
  nor2 g12567(.a(new_n12481), .b(new_n12474), .O(new_n12761));
  nor2 g12568(.a(new_n12761), .b(new_n12760), .O(new_n12762));
  inv1 g12569(.a(new_n12761), .O(new_n12763));
  nor2 g12570(.a(new_n12763), .b(new_n12759), .O(new_n12764));
  nor2 g12571(.a(new_n12764), .b(new_n12762), .O(new_n12765));
  inv1 g12572(.a(new_n12765), .O(new_n12766));
  nor2 g12573(.a(new_n10468), .b(new_n257), .O(new_n12767));
  inv1 g12574(.a(new_n12767), .O(new_n12768));
  nor2 g12575(.a(new_n9873), .b(new_n322), .O(new_n12769));
  nor2 g12576(.a(new_n12769), .b(new_n12389), .O(new_n12770));
  inv1 g12577(.a(new_n12387), .O(new_n12771));
  nor2 g12578(.a(new_n10320), .b(new_n322), .O(new_n12772));
  inv1 g12579(.a(new_n12772), .O(new_n12773));
  nor2 g12580(.a(new_n12773), .b(new_n12771), .O(new_n12774));
  nor2 g12581(.a(new_n12774), .b(new_n12770), .O(new_n12775));
  nor2 g12582(.a(new_n12775), .b(new_n12768), .O(new_n12776));
  inv1 g12583(.a(new_n12775), .O(new_n12777));
  nor2 g12584(.a(new_n12777), .b(new_n12767), .O(new_n12778));
  nor2 g12585(.a(new_n12778), .b(new_n12776), .O(new_n12779));
  nor2 g12586(.a(new_n12779), .b(new_n12766), .O(new_n12780));
  inv1 g12587(.a(new_n12779), .O(new_n12781));
  nor2 g12588(.a(new_n12781), .b(new_n12765), .O(new_n12782));
  nor2 g12589(.a(new_n12782), .b(new_n12780), .O(new_n12783));
  inv1 g12590(.a(new_n12783), .O(new_n12784));
  nor2 g12591(.a(new_n12784), .b(new_n12758), .O(new_n12785));
  inv1 g12592(.a(new_n12758), .O(new_n12786));
  nor2 g12593(.a(new_n12783), .b(new_n12786), .O(new_n12787));
  nor2 g12594(.a(new_n12787), .b(new_n12785), .O(new_n12788));
  nor2 g12595(.a(new_n12788), .b(new_n12757), .O(new_n12789));
  inv1 g12596(.a(new_n12788), .O(new_n12790));
  nor2 g12597(.a(new_n12790), .b(new_n12756), .O(new_n12791));
  nor2 g12598(.a(new_n12791), .b(new_n12789), .O(new_n12792));
  inv1 g12599(.a(new_n12792), .O(new_n12793));
  nor2 g12600(.a(new_n12459), .b(new_n12455), .O(new_n12794));
  nor2 g12601(.a(new_n12443), .b(new_n12435), .O(new_n12795));
  nor2 g12602(.a(new_n12795), .b(new_n12794), .O(new_n12796));
  inv1 g12603(.a(new_n12794), .O(new_n12797));
  inv1 g12604(.a(new_n12795), .O(new_n12798));
  nor2 g12605(.a(new_n12798), .b(new_n12797), .O(new_n12799));
  nor2 g12606(.a(new_n12799), .b(new_n12796), .O(new_n12800));
  nor2 g12607(.a(new_n12321), .b(new_n12316), .O(new_n12801));
  nor2 g12608(.a(new_n12801), .b(new_n12800), .O(new_n12802));
  inv1 g12609(.a(new_n12800), .O(new_n12803));
  inv1 g12610(.a(new_n12801), .O(new_n12804));
  nor2 g12611(.a(new_n12804), .b(new_n12803), .O(new_n12805));
  nor2 g12612(.a(new_n12805), .b(new_n12802), .O(new_n12806));
  inv1 g12613(.a(new_n12806), .O(new_n12807));
  nor2 g12614(.a(new_n12428), .b(new_n12425), .O(new_n12808));
  inv1 g12615(.a(new_n12808), .O(new_n12809));
  nor2 g12616(.a(new_n12408), .b(new_n12400), .O(new_n12810));
  nor2 g12617(.a(new_n12395), .b(new_n12388), .O(new_n12811));
  nor2 g12618(.a(new_n12811), .b(new_n12810), .O(new_n12812));
  inv1 g12619(.a(new_n12810), .O(new_n12813));
  inv1 g12620(.a(new_n12811), .O(new_n12814));
  nor2 g12621(.a(new_n12814), .b(new_n12813), .O(new_n12815));
  nor2 g12622(.a(new_n12815), .b(new_n12812), .O(new_n12816));
  nor2 g12623(.a(new_n12816), .b(new_n12809), .O(new_n12817));
  inv1 g12624(.a(new_n12816), .O(new_n12818));
  nor2 g12625(.a(new_n12818), .b(new_n12808), .O(new_n12819));
  nor2 g12626(.a(new_n12819), .b(new_n12817), .O(new_n12820));
  nor2 g12627(.a(new_n12461), .b(new_n12445), .O(new_n12821));
  inv1 g12628(.a(new_n12821), .O(new_n12822));
  nor2 g12629(.a(new_n12822), .b(new_n12820), .O(new_n12823));
  inv1 g12630(.a(new_n12820), .O(new_n12824));
  nor2 g12631(.a(new_n12821), .b(new_n12824), .O(new_n12825));
  nor2 g12632(.a(new_n12825), .b(new_n12823), .O(new_n12826));
  inv1 g12633(.a(new_n12826), .O(new_n12827));
  nor2 g12634(.a(new_n12827), .b(new_n12807), .O(new_n12828));
  nor2 g12635(.a(new_n12826), .b(new_n12806), .O(new_n12829));
  nor2 g12636(.a(new_n12829), .b(new_n12828), .O(new_n12830));
  inv1 g12637(.a(new_n12830), .O(new_n12831));
  nor2 g12638(.a(new_n12831), .b(new_n12793), .O(new_n12832));
  nor2 g12639(.a(new_n12830), .b(new_n12792), .O(new_n12833));
  nor2 g12640(.a(new_n12833), .b(new_n12832), .O(new_n12834));
  inv1 g12641(.a(new_n12834), .O(new_n12835));
  nor2 g12642(.a(new_n12835), .b(new_n12755), .O(new_n12836));
  inv1 g12643(.a(new_n12755), .O(new_n12837));
  nor2 g12644(.a(new_n12834), .b(new_n12837), .O(new_n12838));
  nor2 g12645(.a(new_n12838), .b(new_n12836), .O(new_n12839));
  inv1 g12646(.a(new_n12839), .O(new_n12840));
  nor2 g12647(.a(new_n12348), .b(new_n12288), .O(new_n12841));
  nor2 g12648(.a(new_n12332), .b(new_n12325), .O(new_n12842));
  nor2 g12649(.a(new_n12508), .b(new_n12501), .O(new_n12843));
  nor2 g12650(.a(new_n12843), .b(new_n12842), .O(new_n12844));
  inv1 g12651(.a(new_n12842), .O(new_n12845));
  inv1 g12652(.a(new_n12843), .O(new_n12846));
  nor2 g12653(.a(new_n12846), .b(new_n12845), .O(new_n12847));
  nor2 g12654(.a(new_n12847), .b(new_n12844), .O(new_n12848));
  nor2 g12655(.a(new_n12495), .b(new_n12487), .O(new_n12849));
  nor2 g12656(.a(new_n12849), .b(new_n12848), .O(new_n12850));
  inv1 g12657(.a(new_n12848), .O(new_n12851));
  inv1 g12658(.a(new_n12849), .O(new_n12852));
  nor2 g12659(.a(new_n12852), .b(new_n12851), .O(new_n12853));
  nor2 g12660(.a(new_n12853), .b(new_n12850), .O(new_n12854));
  nor2 g12661(.a(new_n12417), .b(new_n12411), .O(new_n12855));
  inv1 g12662(.a(new_n12855), .O(new_n12856));
  nor2 g12663(.a(new_n12856), .b(new_n12854), .O(new_n12857));
  inv1 g12664(.a(new_n12854), .O(new_n12858));
  nor2 g12665(.a(new_n12855), .b(new_n12858), .O(new_n12859));
  nor2 g12666(.a(new_n12859), .b(new_n12857), .O(new_n12860));
  nor2 g12667(.a(new_n12517), .b(new_n12510), .O(new_n12861));
  inv1 g12668(.a(new_n12861), .O(new_n12862));
  nor2 g12669(.a(new_n12862), .b(new_n12860), .O(new_n12863));
  inv1 g12670(.a(new_n12860), .O(new_n12864));
  nor2 g12671(.a(new_n12861), .b(new_n12864), .O(new_n12865));
  nor2 g12672(.a(new_n12865), .b(new_n12863), .O(new_n12866));
  inv1 g12673(.a(new_n12866), .O(new_n12867));
  nor2 g12674(.a(new_n12344), .b(new_n12298), .O(new_n12868));
  inv1 g12675(.a(new_n12868), .O(new_n12869));
  nor2 g12676(.a(new_n12520), .b(new_n12466), .O(new_n12870));
  inv1 g12677(.a(new_n12870), .O(new_n12871));
  nor2 g12678(.a(new_n12871), .b(new_n12869), .O(new_n12872));
  nor2 g12679(.a(new_n12870), .b(new_n12868), .O(new_n12873));
  nor2 g12680(.a(new_n12873), .b(new_n12872), .O(new_n12874));
  inv1 g12681(.a(new_n12874), .O(new_n12875));
  nor2 g12682(.a(new_n12875), .b(new_n12867), .O(new_n12876));
  nor2 g12683(.a(new_n12874), .b(new_n12866), .O(new_n12877));
  nor2 g12684(.a(new_n12877), .b(new_n12876), .O(new_n12878));
  inv1 g12685(.a(new_n12878), .O(new_n12879));
  nor2 g12686(.a(new_n12879), .b(new_n12841), .O(new_n12880));
  inv1 g12687(.a(new_n12841), .O(new_n12881));
  nor2 g12688(.a(new_n12878), .b(new_n12881), .O(new_n12882));
  nor2 g12689(.a(new_n12882), .b(new_n12880), .O(new_n12883));
  inv1 g12690(.a(new_n12883), .O(new_n12884));
  nor2 g12691(.a(new_n12884), .b(new_n12840), .O(new_n12885));
  nor2 g12692(.a(new_n12883), .b(new_n12839), .O(new_n12886));
  nor2 g12693(.a(new_n12886), .b(new_n12885), .O(new_n12887));
  inv1 g12694(.a(new_n12887), .O(new_n12888));
  nor2 g12695(.a(new_n12888), .b(new_n12754), .O(new_n12889));
  inv1 g12696(.a(new_n12754), .O(new_n12890));
  nor2 g12697(.a(new_n12887), .b(new_n12890), .O(new_n12891));
  nor2 g12698(.a(new_n12891), .b(new_n12889), .O(new_n12892));
  inv1 g12699(.a(new_n12892), .O(new_n12893));
  nor2 g12700(.a(new_n12893), .b(new_n12753), .O(new_n12894));
  nor2 g12701(.a(new_n12892), .b(new_n12752), .O(new_n12895));
  nor2 g12702(.a(new_n12895), .b(new_n12894), .O(new_n12896));
  inv1 g12703(.a(new_n12896), .O(new_n12897));
  nor2 g12704(.a(new_n12897), .b(new_n12552), .O(new_n12898));
  inv1 g12705(.a(new_n12552), .O(new_n12899));
  nor2 g12706(.a(new_n12896), .b(new_n12899), .O(new_n12900));
  nor2 g12707(.a(new_n12900), .b(new_n12898), .O(new_n12901));
  nor2 g12708(.a(new_n12547), .b(new_n12543), .O(new_n12902));
  inv1 g12709(.a(new_n12902), .O(new_n12903));
  nor2 g12710(.a(new_n12903), .b(new_n12901), .O(new_n12904));
  inv1 g12711(.a(new_n12901), .O(new_n12905));
  nor2 g12712(.a(new_n12902), .b(new_n12905), .O(new_n12906));
  nor2 g12713(.a(new_n12906), .b(new_n12904), .O(new_n12907));
  inv1 g12714(.a(new_n12907), .O(\asquared[67] ));
  nor2 g12715(.a(new_n12894), .b(new_n12889), .O(new_n12909));
  nor2 g12716(.a(new_n12750), .b(new_n12558), .O(new_n12910));
  nor2 g12717(.a(new_n12836), .b(new_n12832), .O(new_n12911));
  inv1 g12718(.a(new_n12911), .O(new_n12912));
  nor2 g12719(.a(new_n12742), .b(new_n12736), .O(new_n12913));
  nor2 g12720(.a(new_n12608), .b(new_n12601), .O(new_n12914));
  inv1 g12721(.a(new_n12914), .O(new_n12915));
  nor2 g12722(.a(new_n12780), .b(new_n12764), .O(new_n12916));
  inv1 g12723(.a(new_n12916), .O(new_n12917));
  nor2 g12724(.a(new_n12917), .b(new_n12915), .O(new_n12918));
  nor2 g12725(.a(new_n12916), .b(new_n12914), .O(new_n12919));
  nor2 g12726(.a(new_n12919), .b(new_n12918), .O(new_n12920));
  nor2 g12727(.a(new_n12708), .b(new_n12701), .O(new_n12921));
  inv1 g12728(.a(new_n12921), .O(new_n12922));
  nor2 g12729(.a(new_n12922), .b(new_n12920), .O(new_n12923));
  inv1 g12730(.a(new_n12920), .O(new_n12924));
  nor2 g12731(.a(new_n12921), .b(new_n12924), .O(new_n12925));
  nor2 g12732(.a(new_n12925), .b(new_n12923), .O(new_n12926));
  inv1 g12733(.a(new_n12926), .O(new_n12927));
  nor2 g12734(.a(new_n12778), .b(new_n12770), .O(new_n12928));
  nor2 g12735(.a(new_n12684), .b(new_n12678), .O(new_n12929));
  nor2 g12736(.a(new_n12929), .b(new_n12928), .O(new_n12930));
  inv1 g12737(.a(new_n12928), .O(new_n12931));
  inv1 g12738(.a(new_n12929), .O(new_n12932));
  nor2 g12739(.a(new_n12932), .b(new_n12931), .O(new_n12933));
  nor2 g12740(.a(new_n12933), .b(new_n12930), .O(new_n12934));
  nor2 g12741(.a(new_n12699), .b(new_n12691), .O(new_n12935));
  nor2 g12742(.a(new_n12935), .b(new_n12934), .O(new_n12936));
  inv1 g12743(.a(new_n12934), .O(new_n12937));
  inv1 g12744(.a(new_n12935), .O(new_n12938));
  nor2 g12745(.a(new_n12938), .b(new_n12937), .O(new_n12939));
  nor2 g12746(.a(new_n12939), .b(new_n12936), .O(new_n12940));
  inv1 g12747(.a(new_n12940), .O(new_n12941));
  nor2 g12748(.a(new_n12572), .b(new_n12565), .O(new_n12942));
  nor2 g12749(.a(new_n12584), .b(new_n12578), .O(new_n12943));
  nor2 g12750(.a(new_n12943), .b(new_n12942), .O(new_n12944));
  inv1 g12751(.a(new_n12942), .O(new_n12945));
  inv1 g12752(.a(new_n12943), .O(new_n12946));
  nor2 g12753(.a(new_n12946), .b(new_n12945), .O(new_n12947));
  nor2 g12754(.a(new_n12947), .b(new_n12944), .O(new_n12948));
  nor2 g12755(.a(new_n12599), .b(new_n12591), .O(new_n12949));
  nor2 g12756(.a(new_n12949), .b(new_n12948), .O(new_n12950));
  inv1 g12757(.a(new_n12948), .O(new_n12951));
  inv1 g12758(.a(new_n12949), .O(new_n12952));
  nor2 g12759(.a(new_n12952), .b(new_n12951), .O(new_n12953));
  nor2 g12760(.a(new_n12953), .b(new_n12950), .O(new_n12954));
  inv1 g12761(.a(new_n12954), .O(new_n12955));
  nor2 g12762(.a(new_n10895), .b(new_n257), .O(new_n12956));
  inv1 g12763(.a(new_n12956), .O(new_n12957));
  nor2 g12764(.a(new_n12619), .b(new_n12612), .O(new_n12958));
  inv1 g12765(.a(new_n12958), .O(new_n12959));
  nor2 g12766(.a(new_n12959), .b(new_n12957), .O(new_n12960));
  nor2 g12767(.a(new_n12958), .b(new_n12956), .O(new_n12961));
  nor2 g12768(.a(new_n12961), .b(new_n12960), .O(new_n12962));
  nor2 g12769(.a(new_n12645), .b(new_n12638), .O(new_n12963));
  nor2 g12770(.a(new_n12963), .b(new_n12962), .O(new_n12964));
  inv1 g12771(.a(new_n12962), .O(new_n12965));
  inv1 g12772(.a(new_n12963), .O(new_n12966));
  nor2 g12773(.a(new_n12966), .b(new_n12965), .O(new_n12967));
  nor2 g12774(.a(new_n12967), .b(new_n12964), .O(new_n12968));
  inv1 g12775(.a(new_n12968), .O(new_n12969));
  nor2 g12776(.a(new_n12969), .b(new_n12955), .O(new_n12970));
  nor2 g12777(.a(new_n12968), .b(new_n12954), .O(new_n12971));
  nor2 g12778(.a(new_n12971), .b(new_n12970), .O(new_n12972));
  inv1 g12779(.a(new_n12972), .O(new_n12973));
  nor2 g12780(.a(new_n12973), .b(new_n12941), .O(new_n12974));
  nor2 g12781(.a(new_n12972), .b(new_n12940), .O(new_n12975));
  nor2 g12782(.a(new_n12975), .b(new_n12974), .O(new_n12976));
  inv1 g12783(.a(new_n12976), .O(new_n12977));
  nor2 g12784(.a(new_n12977), .b(new_n12927), .O(new_n12978));
  nor2 g12785(.a(new_n12976), .b(new_n12926), .O(new_n12979));
  nor2 g12786(.a(new_n12979), .b(new_n12978), .O(new_n12980));
  inv1 g12787(.a(new_n12980), .O(new_n12981));
  nor2 g12788(.a(new_n12981), .b(new_n12913), .O(new_n12982));
  inv1 g12789(.a(new_n12913), .O(new_n12983));
  nor2 g12790(.a(new_n12980), .b(new_n12983), .O(new_n12984));
  nor2 g12791(.a(new_n12984), .b(new_n12982), .O(new_n12985));
  nor2 g12792(.a(new_n12985), .b(new_n12912), .O(new_n12986));
  inv1 g12793(.a(new_n12985), .O(new_n12987));
  nor2 g12794(.a(new_n12987), .b(new_n12911), .O(new_n12988));
  nor2 g12795(.a(new_n12988), .b(new_n12986), .O(new_n12989));
  inv1 g12796(.a(new_n12989), .O(new_n12990));
  nor2 g12797(.a(new_n12672), .b(new_n12665), .O(new_n12991));
  nor2 g12798(.a(new_n12630), .b(new_n12624), .O(new_n12992));
  nor2 g12799(.a(new_n12992), .b(new_n12991), .O(new_n12993));
  inv1 g12800(.a(new_n12991), .O(new_n12994));
  inv1 g12801(.a(new_n12992), .O(new_n12995));
  nor2 g12802(.a(new_n12995), .b(new_n12994), .O(new_n12996));
  nor2 g12803(.a(new_n12996), .b(new_n12993), .O(new_n12997));
  inv1 g12804(.a(new_n12997), .O(new_n12998));
  nor2 g12805(.a(new_n9658), .b(new_n438), .O(new_n12999));
  inv1 g12806(.a(new_n12999), .O(new_n13000));
  nor2 g12807(.a(new_n9156), .b(new_n502), .O(new_n13001));
  nor2 g12808(.a(new_n6570), .b(new_n1297), .O(new_n13002));
  nor2 g12809(.a(new_n13002), .b(new_n13001), .O(new_n13003));
  nor2 g12810(.a(new_n9156), .b(new_n1297), .O(new_n13004));
  inv1 g12811(.a(new_n13004), .O(new_n13005));
  nor2 g12812(.a(new_n13005), .b(new_n11236), .O(new_n13006));
  nor2 g12813(.a(new_n13006), .b(new_n13003), .O(new_n13007));
  nor2 g12814(.a(new_n13007), .b(new_n13000), .O(new_n13008));
  inv1 g12815(.a(new_n13007), .O(new_n13009));
  nor2 g12816(.a(new_n13009), .b(new_n12999), .O(new_n13010));
  nor2 g12817(.a(new_n13010), .b(new_n13008), .O(new_n13011));
  inv1 g12818(.a(new_n13011), .O(new_n13012));
  nor2 g12819(.a(new_n13012), .b(new_n12998), .O(new_n13013));
  nor2 g12820(.a(new_n13011), .b(new_n12997), .O(new_n13014));
  nor2 g12821(.a(new_n13014), .b(new_n13013), .O(new_n13015));
  inv1 g12822(.a(new_n13015), .O(new_n13016));
  nor2 g12823(.a(new_n12654), .b(new_n12647), .O(new_n13017));
  inv1 g12824(.a(new_n13017), .O(new_n13018));
  nor2 g12825(.a(new_n13018), .b(new_n13016), .O(new_n13019));
  nor2 g12826(.a(new_n13017), .b(new_n13015), .O(new_n13020));
  nor2 g12827(.a(new_n13020), .b(new_n13019), .O(new_n13021));
  nor2 g12828(.a(new_n12731), .b(new_n12725), .O(new_n13022));
  inv1 g12829(.a(new_n13022), .O(new_n13023));
  nor2 g12830(.a(new_n13023), .b(new_n13021), .O(new_n13024));
  inv1 g12831(.a(new_n13021), .O(new_n13025));
  nor2 g12832(.a(new_n13022), .b(new_n13025), .O(new_n13026));
  nor2 g12833(.a(new_n13026), .b(new_n13024), .O(new_n13027));
  inv1 g12834(.a(new_n13027), .O(new_n13028));
  nor2 g12835(.a(new_n12711), .b(new_n12657), .O(new_n13029));
  inv1 g12836(.a(new_n13029), .O(new_n13030));
  nor2 g12837(.a(new_n12791), .b(new_n12785), .O(new_n13031));
  inv1 g12838(.a(new_n13031), .O(new_n13032));
  nor2 g12839(.a(new_n13032), .b(new_n13030), .O(new_n13033));
  nor2 g12840(.a(new_n13031), .b(new_n13029), .O(new_n13034));
  nor2 g12841(.a(new_n13034), .b(new_n13033), .O(new_n13035));
  inv1 g12842(.a(new_n13035), .O(new_n13036));
  nor2 g12843(.a(new_n13036), .b(new_n13028), .O(new_n13037));
  nor2 g12844(.a(new_n13035), .b(new_n13027), .O(new_n13038));
  nor2 g12845(.a(new_n13038), .b(new_n13037), .O(new_n13039));
  inv1 g12846(.a(new_n13039), .O(new_n13040));
  nor2 g12847(.a(new_n13040), .b(new_n12990), .O(new_n13041));
  nor2 g12848(.a(new_n13039), .b(new_n12989), .O(new_n13042));
  nor2 g12849(.a(new_n13042), .b(new_n13041), .O(new_n13043));
  inv1 g12850(.a(new_n13043), .O(new_n13044));
  nor2 g12851(.a(new_n13044), .b(new_n12910), .O(new_n13045));
  inv1 g12852(.a(new_n12910), .O(new_n13046));
  nor2 g12853(.a(new_n13043), .b(new_n13046), .O(new_n13047));
  nor2 g12854(.a(new_n13047), .b(new_n13045), .O(new_n13048));
  inv1 g12855(.a(new_n13048), .O(new_n13049));
  nor2 g12856(.a(new_n12885), .b(new_n12880), .O(new_n13050));
  inv1 g12857(.a(new_n13050), .O(new_n13051));
  nor2 g12858(.a(new_n12746), .b(new_n12715), .O(new_n13052));
  inv1 g12859(.a(new_n13052), .O(new_n13053));
  nor2 g12860(.a(new_n13053), .b(new_n13051), .O(new_n13054));
  nor2 g12861(.a(new_n13052), .b(new_n13050), .O(new_n13055));
  nor2 g12862(.a(new_n13055), .b(new_n13054), .O(new_n13056));
  inv1 g12863(.a(new_n13056), .O(new_n13057));
  nor2 g12864(.a(new_n12876), .b(new_n12873), .O(new_n13058));
  nor2 g12865(.a(new_n4682), .b(new_n2184), .O(new_n13059));
  nor2 g12866(.a(new_n4425), .b(new_n2433), .O(new_n13060));
  nor2 g12867(.a(new_n13060), .b(new_n13059), .O(new_n13061));
  nor2 g12868(.a(new_n4682), .b(new_n2433), .O(new_n13062));
  inv1 g12869(.a(new_n13062), .O(new_n13063));
  nor2 g12870(.a(new_n13063), .b(new_n12689), .O(new_n13064));
  nor2 g12871(.a(new_n13064), .b(new_n13061), .O(new_n13065));
  nor2 g12872(.a(new_n13065), .b(new_n12304), .O(new_n13066));
  inv1 g12873(.a(new_n13065), .O(new_n13067));
  nor2 g12874(.a(new_n13067), .b(new_n12303), .O(new_n13068));
  nor2 g12875(.a(new_n13068), .b(new_n13066), .O(new_n13069));
  nor2 g12876(.a(new_n5178), .b(new_n1903), .O(new_n13070));
  inv1 g12877(.a(new_n13070), .O(new_n13071));
  nor2 g12878(.a(new_n6274), .b(new_n1425), .O(new_n13072));
  nor2 g12879(.a(new_n13072), .b(new_n12566), .O(new_n13073));
  inv1 g12880(.a(new_n13072), .O(new_n13074));
  nor2 g12881(.a(new_n13074), .b(new_n12567), .O(new_n13075));
  nor2 g12882(.a(new_n13075), .b(new_n13073), .O(new_n13076));
  nor2 g12883(.a(new_n13076), .b(new_n13071), .O(new_n13077));
  inv1 g12884(.a(new_n13076), .O(new_n13078));
  nor2 g12885(.a(new_n13078), .b(new_n13070), .O(new_n13079));
  nor2 g12886(.a(new_n13079), .b(new_n13077), .O(new_n13080));
  nor2 g12887(.a(new_n6893), .b(new_n1199), .O(new_n13081));
  inv1 g12888(.a(new_n13081), .O(new_n13082));
  nor2 g12889(.a(new_n8170), .b(new_n699), .O(new_n13083));
  nor2 g12890(.a(new_n13083), .b(new_n12613), .O(new_n13084));
  inv1 g12891(.a(new_n13083), .O(new_n13085));
  nor2 g12892(.a(new_n13085), .b(new_n12614), .O(new_n13086));
  nor2 g12893(.a(new_n13086), .b(new_n13084), .O(new_n13087));
  nor2 g12894(.a(new_n13087), .b(new_n13082), .O(new_n13088));
  inv1 g12895(.a(new_n13087), .O(new_n13089));
  nor2 g12896(.a(new_n13089), .b(new_n13081), .O(new_n13090));
  nor2 g12897(.a(new_n13090), .b(new_n13088), .O(new_n13091));
  nor2 g12898(.a(new_n13091), .b(new_n13080), .O(new_n13092));
  inv1 g12899(.a(new_n13080), .O(new_n13093));
  inv1 g12900(.a(new_n13091), .O(new_n13094));
  nor2 g12901(.a(new_n13094), .b(new_n13093), .O(new_n13095));
  nor2 g12902(.a(new_n13095), .b(new_n13092), .O(new_n13096));
  inv1 g12903(.a(new_n13096), .O(new_n13097));
  nor2 g12904(.a(new_n13097), .b(new_n13069), .O(new_n13098));
  inv1 g12905(.a(new_n13069), .O(new_n13099));
  nor2 g12906(.a(new_n13096), .b(new_n13099), .O(new_n13100));
  nor2 g12907(.a(new_n13100), .b(new_n13098), .O(new_n13101));
  inv1 g12908(.a(new_n13101), .O(new_n13102));
  nor2 g12909(.a(new_n8946), .b(new_n569), .O(new_n13103));
  nor2 g12910(.a(new_n8476), .b(new_n613), .O(new_n13104));
  nor2 g12911(.a(new_n13104), .b(new_n13103), .O(new_n13105));
  nor2 g12912(.a(new_n8946), .b(new_n613), .O(new_n13106));
  inv1 g12913(.a(new_n13106), .O(new_n13107));
  nor2 g12914(.a(new_n13107), .b(new_n12667), .O(new_n13108));
  nor2 g12915(.a(new_n13108), .b(new_n13105), .O(new_n13109));
  nor2 g12916(.a(new_n13109), .b(new_n12694), .O(new_n13110));
  inv1 g12917(.a(new_n13109), .O(new_n13111));
  nor2 g12918(.a(new_n13111), .b(new_n12693), .O(new_n13112));
  nor2 g12919(.a(new_n13112), .b(new_n13110), .O(new_n13113));
  nor2 g12920(.a(new_n3533), .b(new_n3231), .O(new_n13114));
  nor2 g12921(.a(new_n3722), .b(new_n3057), .O(new_n13115));
  nor2 g12922(.a(new_n13115), .b(new_n13114), .O(new_n13116));
  nor2 g12923(.a(new_n3722), .b(new_n3231), .O(new_n13117));
  inv1 g12924(.a(new_n13117), .O(new_n13118));
  nor2 g12925(.a(new_n13118), .b(new_n12438), .O(new_n13119));
  nor2 g12926(.a(new_n13119), .b(new_n13116), .O(new_n13120));
  nor2 g12927(.a(new_n13120), .b(new_n12640), .O(new_n13121));
  inv1 g12928(.a(new_n13120), .O(new_n13122));
  nor2 g12929(.a(new_n13122), .b(new_n12639), .O(new_n13123));
  nor2 g12930(.a(new_n13123), .b(new_n13121), .O(new_n13124));
  nor2 g12931(.a(new_n6958), .b(new_n1086), .O(new_n13125));
  inv1 g12932(.a(new_n13125), .O(new_n13126));
  nor2 g12933(.a(new_n12679), .b(\a[34] ), .O(new_n13127));
  inv1 g12934(.a(new_n4604), .O(new_n13128));
  nor2 g12935(.a(new_n13128), .b(new_n11186), .O(new_n13129));
  nor2 g12936(.a(new_n13129), .b(new_n13127), .O(new_n13130));
  nor2 g12937(.a(new_n13130), .b(new_n13126), .O(new_n13131));
  nor2 g12938(.a(new_n13127), .b(new_n13126), .O(new_n13132));
  nor2 g12939(.a(new_n13132), .b(new_n13129), .O(new_n13133));
  inv1 g12940(.a(new_n13133), .O(new_n13134));
  nor2 g12941(.a(new_n13134), .b(new_n13127), .O(new_n13135));
  nor2 g12942(.a(new_n13135), .b(new_n13131), .O(new_n13136));
  nor2 g12943(.a(new_n13136), .b(new_n13124), .O(new_n13137));
  inv1 g12944(.a(new_n13124), .O(new_n13138));
  inv1 g12945(.a(new_n13136), .O(new_n13139));
  nor2 g12946(.a(new_n13139), .b(new_n13138), .O(new_n13140));
  nor2 g12947(.a(new_n13140), .b(new_n13137), .O(new_n13141));
  inv1 g12948(.a(new_n13141), .O(new_n13142));
  nor2 g12949(.a(new_n13142), .b(new_n13113), .O(new_n13143));
  inv1 g12950(.a(new_n13113), .O(new_n13144));
  nor2 g12951(.a(new_n13141), .b(new_n13144), .O(new_n13145));
  nor2 g12952(.a(new_n13145), .b(new_n13143), .O(new_n13146));
  inv1 g12953(.a(new_n13146), .O(new_n13147));
  nor2 g12954(.a(new_n8026), .b(new_n800), .O(new_n13148));
  inv1 g12955(.a(new_n13148), .O(new_n13149));
  nor2 g12956(.a(new_n4093), .b(new_n2660), .O(new_n13150));
  nor2 g12957(.a(new_n13150), .b(new_n10615), .O(new_n13151));
  inv1 g12958(.a(new_n13150), .O(new_n13152));
  nor2 g12959(.a(new_n13152), .b(new_n10616), .O(new_n13153));
  nor2 g12960(.a(new_n13153), .b(new_n13151), .O(new_n13154));
  nor2 g12961(.a(new_n13154), .b(new_n13149), .O(new_n13155));
  inv1 g12962(.a(new_n13154), .O(new_n13156));
  nor2 g12963(.a(new_n13156), .b(new_n13148), .O(new_n13157));
  nor2 g12964(.a(new_n13157), .b(new_n13155), .O(new_n13158));
  inv1 g12965(.a(new_n13158), .O(new_n13159));
  nor2 g12966(.a(new_n10468), .b(new_n295), .O(new_n13160));
  nor2 g12967(.a(new_n9873), .b(new_n363), .O(new_n13161));
  nor2 g12968(.a(new_n13161), .b(new_n12772), .O(new_n13162));
  inv1 g12969(.a(new_n12769), .O(new_n13163));
  nor2 g12970(.a(new_n10320), .b(new_n363), .O(new_n13164));
  inv1 g12971(.a(new_n13164), .O(new_n13165));
  nor2 g12972(.a(new_n13165), .b(new_n13163), .O(new_n13166));
  nor2 g12973(.a(new_n13166), .b(new_n13162), .O(new_n13167));
  inv1 g12974(.a(new_n13167), .O(new_n13168));
  nor2 g12975(.a(new_n13168), .b(new_n13160), .O(new_n13169));
  inv1 g12976(.a(new_n13160), .O(new_n13170));
  nor2 g12977(.a(new_n13167), .b(new_n13170), .O(new_n13171));
  nor2 g12978(.a(new_n13171), .b(new_n13169), .O(new_n13172));
  nor2 g12979(.a(new_n5796), .b(new_n1647), .O(new_n13173));
  nor2 g12980(.a(new_n5393), .b(new_n1736), .O(new_n13174));
  nor2 g12981(.a(new_n13174), .b(new_n13173), .O(new_n13175));
  nor2 g12982(.a(new_n5796), .b(new_n1736), .O(new_n13176));
  inv1 g12983(.a(new_n13176), .O(new_n13177));
  nor2 g12984(.a(new_n13177), .b(new_n12585), .O(new_n13178));
  nor2 g12985(.a(new_n13178), .b(new_n13175), .O(new_n13179));
  nor2 g12986(.a(new_n13179), .b(new_n12594), .O(new_n13180));
  inv1 g12987(.a(new_n13179), .O(new_n13181));
  nor2 g12988(.a(new_n13181), .b(new_n12593), .O(new_n13182));
  nor2 g12989(.a(new_n13182), .b(new_n13180), .O(new_n13183));
  nor2 g12990(.a(new_n13183), .b(new_n13172), .O(new_n13184));
  inv1 g12991(.a(new_n13172), .O(new_n13185));
  inv1 g12992(.a(new_n13183), .O(new_n13186));
  nor2 g12993(.a(new_n13186), .b(new_n13185), .O(new_n13187));
  nor2 g12994(.a(new_n13187), .b(new_n13184), .O(new_n13188));
  nor2 g12995(.a(new_n13188), .b(new_n13159), .O(new_n13189));
  inv1 g12996(.a(new_n13188), .O(new_n13190));
  nor2 g12997(.a(new_n13190), .b(new_n13158), .O(new_n13191));
  nor2 g12998(.a(new_n13191), .b(new_n13189), .O(new_n13192));
  inv1 g12999(.a(new_n13192), .O(new_n13193));
  nor2 g13000(.a(new_n13193), .b(new_n13147), .O(new_n13194));
  nor2 g13001(.a(new_n13192), .b(new_n13146), .O(new_n13195));
  nor2 g13002(.a(new_n13195), .b(new_n13194), .O(new_n13196));
  inv1 g13003(.a(new_n13196), .O(new_n13197));
  nor2 g13004(.a(new_n13197), .b(new_n13102), .O(new_n13198));
  nor2 g13005(.a(new_n13196), .b(new_n13101), .O(new_n13199));
  nor2 g13006(.a(new_n13199), .b(new_n13198), .O(new_n13200));
  inv1 g13007(.a(new_n13200), .O(new_n13201));
  nor2 g13008(.a(new_n13201), .b(new_n13058), .O(new_n13202));
  inv1 g13009(.a(new_n13058), .O(new_n13203));
  nor2 g13010(.a(new_n13200), .b(new_n13203), .O(new_n13204));
  nor2 g13011(.a(new_n13204), .b(new_n13202), .O(new_n13205));
  inv1 g13012(.a(new_n13205), .O(new_n13206));
  nor2 g13013(.a(new_n12819), .b(new_n12815), .O(new_n13207));
  inv1 g13014(.a(new_n13207), .O(new_n13208));
  nor2 g13015(.a(new_n12853), .b(new_n12847), .O(new_n13209));
  inv1 g13016(.a(new_n13209), .O(new_n13210));
  nor2 g13017(.a(new_n13210), .b(new_n13208), .O(new_n13211));
  nor2 g13018(.a(new_n13209), .b(new_n13207), .O(new_n13212));
  nor2 g13019(.a(new_n13212), .b(new_n13211), .O(new_n13213));
  nor2 g13020(.a(new_n12805), .b(new_n12799), .O(new_n13214));
  inv1 g13021(.a(new_n13214), .O(new_n13215));
  nor2 g13022(.a(new_n13215), .b(new_n13213), .O(new_n13216));
  inv1 g13023(.a(new_n13213), .O(new_n13217));
  nor2 g13024(.a(new_n13214), .b(new_n13217), .O(new_n13218));
  nor2 g13025(.a(new_n13218), .b(new_n13216), .O(new_n13219));
  inv1 g13026(.a(new_n13219), .O(new_n13220));
  nor2 g13027(.a(new_n12828), .b(new_n12825), .O(new_n13221));
  inv1 g13028(.a(new_n13221), .O(new_n13222));
  nor2 g13029(.a(new_n12865), .b(new_n12859), .O(new_n13223));
  inv1 g13030(.a(new_n13223), .O(new_n13224));
  nor2 g13031(.a(new_n13224), .b(new_n13222), .O(new_n13225));
  nor2 g13032(.a(new_n13223), .b(new_n13221), .O(new_n13226));
  nor2 g13033(.a(new_n13226), .b(new_n13225), .O(new_n13227));
  inv1 g13034(.a(new_n13227), .O(new_n13228));
  nor2 g13035(.a(new_n13228), .b(new_n13220), .O(new_n13229));
  nor2 g13036(.a(new_n13227), .b(new_n13219), .O(new_n13230));
  nor2 g13037(.a(new_n13230), .b(new_n13229), .O(new_n13231));
  inv1 g13038(.a(new_n13231), .O(new_n13232));
  nor2 g13039(.a(new_n13232), .b(new_n13206), .O(new_n13233));
  nor2 g13040(.a(new_n13231), .b(new_n13205), .O(new_n13234));
  nor2 g13041(.a(new_n13234), .b(new_n13233), .O(new_n13235));
  inv1 g13042(.a(new_n13235), .O(new_n13236));
  nor2 g13043(.a(new_n13236), .b(new_n13057), .O(new_n13237));
  nor2 g13044(.a(new_n13235), .b(new_n13056), .O(new_n13238));
  nor2 g13045(.a(new_n13238), .b(new_n13237), .O(new_n13239));
  inv1 g13046(.a(new_n13239), .O(new_n13240));
  nor2 g13047(.a(new_n13240), .b(new_n13049), .O(new_n13241));
  nor2 g13048(.a(new_n13239), .b(new_n13048), .O(new_n13242));
  nor2 g13049(.a(new_n13242), .b(new_n13241), .O(new_n13243));
  inv1 g13050(.a(new_n13243), .O(new_n13244));
  nor2 g13051(.a(new_n13244), .b(new_n12909), .O(new_n13245));
  inv1 g13052(.a(new_n12909), .O(new_n13246));
  nor2 g13053(.a(new_n13243), .b(new_n13246), .O(new_n13247));
  nor2 g13054(.a(new_n13247), .b(new_n13245), .O(new_n13248));
  inv1 g13055(.a(new_n13248), .O(new_n13249));
  nor2 g13056(.a(new_n12906), .b(new_n12900), .O(new_n13250));
  nor2 g13057(.a(new_n13250), .b(new_n13249), .O(new_n13251));
  inv1 g13058(.a(new_n13250), .O(new_n13252));
  nor2 g13059(.a(new_n13252), .b(new_n13248), .O(new_n13253));
  nor2 g13060(.a(new_n13253), .b(new_n13251), .O(new_n13254));
  inv1 g13061(.a(new_n13254), .O(\asquared[68] ));
  nor2 g13062(.a(new_n13241), .b(new_n13045), .O(new_n13256));
  inv1 g13063(.a(new_n13256), .O(new_n13257));
  nor2 g13064(.a(new_n13041), .b(new_n12988), .O(new_n13258));
  nor2 g13065(.a(new_n13233), .b(new_n13202), .O(new_n13259));
  nor2 g13066(.a(new_n13037), .b(new_n13034), .O(new_n13260));
  nor2 g13067(.a(new_n12974), .b(new_n12970), .O(new_n13261));
  inv1 g13068(.a(new_n13261), .O(new_n13262));
  nor2 g13069(.a(new_n12925), .b(new_n12919), .O(new_n13263));
  inv1 g13070(.a(new_n13263), .O(new_n13264));
  nor2 g13071(.a(new_n13264), .b(new_n13262), .O(new_n13265));
  nor2 g13072(.a(new_n13263), .b(new_n13261), .O(new_n13266));
  nor2 g13073(.a(new_n13266), .b(new_n13265), .O(new_n13267));
  nor2 g13074(.a(new_n13026), .b(new_n13020), .O(new_n13268));
  inv1 g13075(.a(new_n13268), .O(new_n13269));
  nor2 g13076(.a(new_n13269), .b(new_n13267), .O(new_n13270));
  inv1 g13077(.a(new_n13267), .O(new_n13271));
  nor2 g13078(.a(new_n13268), .b(new_n13271), .O(new_n13272));
  nor2 g13079(.a(new_n13272), .b(new_n13270), .O(new_n13273));
  inv1 g13080(.a(new_n13273), .O(new_n13274));
  nor2 g13081(.a(new_n7294), .b(new_n1086), .O(new_n13275));
  nor2 g13082(.a(new_n6958), .b(new_n1199), .O(new_n13276));
  nor2 g13083(.a(new_n13276), .b(new_n13275), .O(new_n13277));
  nor2 g13084(.a(new_n7294), .b(new_n1199), .O(new_n13278));
  inv1 g13085(.a(new_n13278), .O(new_n13279));
  nor2 g13086(.a(new_n13279), .b(new_n13126), .O(new_n13280));
  nor2 g13087(.a(new_n13280), .b(new_n13277), .O(new_n13281));
  inv1 g13088(.a(new_n13281), .O(new_n13282));
  nor2 g13089(.a(new_n13282), .b(new_n13117), .O(new_n13283));
  nor2 g13090(.a(new_n13281), .b(new_n13118), .O(new_n13284));
  nor2 g13091(.a(new_n13284), .b(new_n13283), .O(new_n13285));
  nor2 g13092(.a(new_n4366), .b(new_n2660), .O(new_n13286));
  inv1 g13093(.a(new_n13286), .O(new_n13287));
  nor2 g13094(.a(new_n3870), .b(new_n3057), .O(new_n13288));
  nor2 g13095(.a(new_n4093), .b(new_n2826), .O(new_n13289));
  nor2 g13096(.a(new_n13289), .b(new_n13288), .O(new_n13290));
  nor2 g13097(.a(new_n4093), .b(new_n3057), .O(new_n13291));
  inv1 g13098(.a(new_n13291), .O(new_n13292));
  nor2 g13099(.a(new_n13292), .b(new_n12640), .O(new_n13293));
  nor2 g13100(.a(new_n13293), .b(new_n13290), .O(new_n13294));
  nor2 g13101(.a(new_n13294), .b(new_n13287), .O(new_n13295));
  inv1 g13102(.a(new_n13294), .O(new_n13296));
  nor2 g13103(.a(new_n13296), .b(new_n13286), .O(new_n13297));
  nor2 g13104(.a(new_n13297), .b(new_n13295), .O(new_n13298));
  nor2 g13105(.a(new_n13298), .b(new_n13285), .O(new_n13299));
  inv1 g13106(.a(new_n13285), .O(new_n13300));
  inv1 g13107(.a(new_n13298), .O(new_n13301));
  nor2 g13108(.a(new_n13301), .b(new_n13300), .O(new_n13302));
  nor2 g13109(.a(new_n13302), .b(new_n13299), .O(new_n13303));
  inv1 g13110(.a(new_n13303), .O(new_n13304));
  nor2 g13111(.a(new_n9156), .b(new_n569), .O(new_n13305));
  inv1 g13112(.a(new_n13305), .O(new_n13306));
  nor2 g13113(.a(new_n13106), .b(new_n9505), .O(new_n13307));
  nor2 g13114(.a(new_n13107), .b(new_n9506), .O(new_n13308));
  nor2 g13115(.a(new_n13308), .b(new_n13307), .O(new_n13309));
  nor2 g13116(.a(new_n13309), .b(new_n13306), .O(new_n13310));
  inv1 g13117(.a(new_n13309), .O(new_n13311));
  nor2 g13118(.a(new_n13311), .b(new_n13305), .O(new_n13312));
  nor2 g13119(.a(new_n13312), .b(new_n13310), .O(new_n13313));
  nor2 g13120(.a(new_n13313), .b(new_n13304), .O(new_n13314));
  inv1 g13121(.a(new_n13313), .O(new_n13315));
  nor2 g13122(.a(new_n13315), .b(new_n13303), .O(new_n13316));
  nor2 g13123(.a(new_n13316), .b(new_n13314), .O(new_n13317));
  inv1 g13124(.a(new_n13317), .O(new_n13318));
  nor2 g13125(.a(new_n5393), .b(new_n1903), .O(new_n13319));
  nor2 g13126(.a(new_n5178), .b(new_n2121), .O(new_n13320));
  nor2 g13127(.a(new_n13320), .b(new_n13319), .O(new_n13321));
  nor2 g13128(.a(new_n5393), .b(new_n2121), .O(new_n13322));
  inv1 g13129(.a(new_n13322), .O(new_n13323));
  nor2 g13130(.a(new_n13323), .b(new_n13071), .O(new_n13324));
  nor2 g13131(.a(new_n13324), .b(new_n13321), .O(new_n13325));
  nor2 g13132(.a(new_n13325), .b(new_n13177), .O(new_n13326));
  inv1 g13133(.a(new_n13325), .O(new_n13327));
  nor2 g13134(.a(new_n13327), .b(new_n13176), .O(new_n13328));
  nor2 g13135(.a(new_n13328), .b(new_n13326), .O(new_n13329));
  inv1 g13136(.a(new_n13329), .O(new_n13330));
  nor2 g13137(.a(new_n8476), .b(new_n699), .O(new_n13331));
  nor2 g13138(.a(new_n12625), .b(new_n11678), .O(new_n13332));
  nor2 g13139(.a(new_n8170), .b(new_n847), .O(new_n13333));
  inv1 g13140(.a(new_n13333), .O(new_n13334));
  nor2 g13141(.a(new_n13334), .b(new_n13149), .O(new_n13335));
  nor2 g13142(.a(new_n13335), .b(new_n13332), .O(new_n13336));
  inv1 g13143(.a(new_n13336), .O(new_n13337));
  nor2 g13144(.a(new_n13337), .b(new_n13331), .O(new_n13338));
  inv1 g13145(.a(new_n13331), .O(new_n13339));
  nor2 g13146(.a(new_n13336), .b(new_n13339), .O(new_n13340));
  nor2 g13147(.a(new_n13340), .b(new_n13338), .O(new_n13341));
  nor2 g13148(.a(new_n6893), .b(new_n1297), .O(new_n13342));
  inv1 g13149(.a(new_n13342), .O(new_n13343));
  nor2 g13150(.a(new_n5971), .b(new_n1647), .O(new_n13344));
  nor2 g13151(.a(new_n6274), .b(new_n1493), .O(new_n13345));
  nor2 g13152(.a(new_n13345), .b(new_n13344), .O(new_n13346));
  nor2 g13153(.a(new_n6274), .b(new_n1647), .O(new_n13347));
  inv1 g13154(.a(new_n13347), .O(new_n13348));
  nor2 g13155(.a(new_n13348), .b(new_n12594), .O(new_n13349));
  nor2 g13156(.a(new_n13349), .b(new_n13346), .O(new_n13350));
  nor2 g13157(.a(new_n13350), .b(new_n13343), .O(new_n13351));
  inv1 g13158(.a(new_n13350), .O(new_n13352));
  nor2 g13159(.a(new_n13352), .b(new_n13342), .O(new_n13353));
  nor2 g13160(.a(new_n13353), .b(new_n13351), .O(new_n13354));
  nor2 g13161(.a(new_n13354), .b(new_n13341), .O(new_n13355));
  inv1 g13162(.a(new_n13341), .O(new_n13356));
  inv1 g13163(.a(new_n13354), .O(new_n13357));
  nor2 g13164(.a(new_n13357), .b(new_n13356), .O(new_n13358));
  nor2 g13165(.a(new_n13358), .b(new_n13355), .O(new_n13359));
  nor2 g13166(.a(new_n13359), .b(new_n13330), .O(new_n13360));
  inv1 g13167(.a(new_n13359), .O(new_n13361));
  nor2 g13168(.a(new_n13361), .b(new_n13329), .O(new_n13362));
  nor2 g13169(.a(new_n13362), .b(new_n13360), .O(new_n13363));
  inv1 g13170(.a(new_n13363), .O(new_n13364));
  nor2 g13171(.a(new_n13364), .b(new_n13318), .O(new_n13365));
  nor2 g13172(.a(new_n13363), .b(new_n13317), .O(new_n13366));
  nor2 g13173(.a(new_n13366), .b(new_n13365), .O(new_n13367));
  inv1 g13174(.a(new_n13367), .O(new_n13368));
  nor2 g13175(.a(new_n6570), .b(new_n1425), .O(new_n13369));
  inv1 g13176(.a(new_n13369), .O(new_n13370));
  nor2 g13177(.a(new_n11596), .b(new_n229), .O(new_n13371));
  nor2 g13178(.a(new_n11186), .b(new_n257), .O(new_n13372));
  nor2 g13179(.a(new_n13372), .b(new_n13371), .O(new_n13373));
  nor2 g13180(.a(new_n11596), .b(new_n257), .O(new_n13374));
  inv1 g13181(.a(new_n13374), .O(new_n13375));
  nor2 g13182(.a(new_n13375), .b(new_n12680), .O(new_n13376));
  nor2 g13183(.a(new_n13376), .b(new_n13373), .O(new_n13377));
  nor2 g13184(.a(new_n13377), .b(new_n13370), .O(new_n13378));
  inv1 g13185(.a(new_n13377), .O(new_n13379));
  nor2 g13186(.a(new_n13379), .b(new_n13369), .O(new_n13380));
  nor2 g13187(.a(new_n13380), .b(new_n13378), .O(new_n13381));
  inv1 g13188(.a(new_n13381), .O(new_n13382));
  nor2 g13189(.a(new_n9873), .b(new_n438), .O(new_n13383));
  nor2 g13190(.a(new_n9658), .b(new_n502), .O(new_n13384));
  nor2 g13191(.a(new_n13384), .b(new_n13383), .O(new_n13385));
  nor2 g13192(.a(new_n9873), .b(new_n502), .O(new_n13386));
  inv1 g13193(.a(new_n13386), .O(new_n13387));
  nor2 g13194(.a(new_n13387), .b(new_n13000), .O(new_n13388));
  nor2 g13195(.a(new_n13388), .b(new_n13385), .O(new_n13389));
  inv1 g13196(.a(new_n13389), .O(new_n13390));
  nor2 g13197(.a(new_n13390), .b(new_n13164), .O(new_n13391));
  nor2 g13198(.a(new_n13389), .b(new_n13165), .O(new_n13392));
  nor2 g13199(.a(new_n13392), .b(new_n13391), .O(new_n13393));
  nor2 g13200(.a(new_n4954), .b(new_n2184), .O(new_n13394));
  inv1 g13201(.a(new_n13394), .O(new_n13395));
  nor2 g13202(.a(new_n4425), .b(new_n2506), .O(new_n13396));
  nor2 g13203(.a(new_n13396), .b(new_n13062), .O(new_n13397));
  inv1 g13204(.a(new_n13060), .O(new_n13398));
  nor2 g13205(.a(new_n4682), .b(new_n2506), .O(new_n13399));
  inv1 g13206(.a(new_n13399), .O(new_n13400));
  nor2 g13207(.a(new_n13400), .b(new_n13398), .O(new_n13401));
  nor2 g13208(.a(new_n13401), .b(new_n13397), .O(new_n13402));
  nor2 g13209(.a(new_n13402), .b(new_n13395), .O(new_n13403));
  inv1 g13210(.a(new_n13402), .O(new_n13404));
  nor2 g13211(.a(new_n13404), .b(new_n13394), .O(new_n13405));
  nor2 g13212(.a(new_n13405), .b(new_n13403), .O(new_n13406));
  nor2 g13213(.a(new_n13406), .b(new_n13393), .O(new_n13407));
  inv1 g13214(.a(new_n13393), .O(new_n13408));
  inv1 g13215(.a(new_n13406), .O(new_n13409));
  nor2 g13216(.a(new_n13409), .b(new_n13408), .O(new_n13410));
  nor2 g13217(.a(new_n13410), .b(new_n13407), .O(new_n13411));
  nor2 g13218(.a(new_n13411), .b(new_n13382), .O(new_n13412));
  inv1 g13219(.a(new_n13411), .O(new_n13413));
  nor2 g13220(.a(new_n13413), .b(new_n13381), .O(new_n13414));
  nor2 g13221(.a(new_n13414), .b(new_n13412), .O(new_n13415));
  inv1 g13222(.a(new_n13415), .O(new_n13416));
  nor2 g13223(.a(new_n13416), .b(new_n13368), .O(new_n13417));
  nor2 g13224(.a(new_n13415), .b(new_n13367), .O(new_n13418));
  nor2 g13225(.a(new_n13418), .b(new_n13417), .O(new_n13419));
  inv1 g13226(.a(new_n13419), .O(new_n13420));
  nor2 g13227(.a(new_n13420), .b(new_n13274), .O(new_n13421));
  nor2 g13228(.a(new_n13419), .b(new_n13273), .O(new_n13422));
  nor2 g13229(.a(new_n13422), .b(new_n13421), .O(new_n13423));
  inv1 g13230(.a(new_n13423), .O(new_n13424));
  nor2 g13231(.a(new_n13424), .b(new_n13260), .O(new_n13425));
  inv1 g13232(.a(new_n13260), .O(new_n13426));
  nor2 g13233(.a(new_n13423), .b(new_n13426), .O(new_n13427));
  nor2 g13234(.a(new_n13427), .b(new_n13425), .O(new_n13428));
  inv1 g13235(.a(new_n13428), .O(new_n13429));
  nor2 g13236(.a(new_n13429), .b(new_n13259), .O(new_n13430));
  inv1 g13237(.a(new_n13259), .O(new_n13431));
  nor2 g13238(.a(new_n13428), .b(new_n13431), .O(new_n13432));
  nor2 g13239(.a(new_n13432), .b(new_n13430), .O(new_n13433));
  inv1 g13240(.a(new_n13433), .O(new_n13434));
  nor2 g13241(.a(new_n13434), .b(new_n13258), .O(new_n13435));
  inv1 g13242(.a(new_n13258), .O(new_n13436));
  nor2 g13243(.a(new_n13433), .b(new_n13436), .O(new_n13437));
  nor2 g13244(.a(new_n13437), .b(new_n13435), .O(new_n13438));
  inv1 g13245(.a(new_n13438), .O(new_n13439));
  nor2 g13246(.a(new_n13237), .b(new_n13055), .O(new_n13440));
  nor2 g13247(.a(new_n13229), .b(new_n13226), .O(new_n13441));
  nor2 g13248(.a(new_n13090), .b(new_n13084), .O(new_n13442));
  nor2 g13249(.a(new_n13079), .b(new_n13073), .O(new_n13443));
  nor2 g13250(.a(new_n13443), .b(new_n13442), .O(new_n13444));
  inv1 g13251(.a(new_n13442), .O(new_n13445));
  inv1 g13252(.a(new_n13443), .O(new_n13446));
  nor2 g13253(.a(new_n13446), .b(new_n13445), .O(new_n13447));
  nor2 g13254(.a(new_n13447), .b(new_n13444), .O(new_n13448));
  nor2 g13255(.a(new_n13112), .b(new_n13105), .O(new_n13449));
  nor2 g13256(.a(new_n13449), .b(new_n13448), .O(new_n13450));
  inv1 g13257(.a(new_n13448), .O(new_n13451));
  inv1 g13258(.a(new_n13449), .O(new_n13452));
  nor2 g13259(.a(new_n13452), .b(new_n13451), .O(new_n13453));
  nor2 g13260(.a(new_n13453), .b(new_n13450), .O(new_n13454));
  inv1 g13261(.a(new_n13454), .O(new_n13455));
  nor2 g13262(.a(new_n13098), .b(new_n13092), .O(new_n13456));
  inv1 g13263(.a(new_n13456), .O(new_n13457));
  nor2 g13264(.a(new_n13143), .b(new_n13137), .O(new_n13458));
  inv1 g13265(.a(new_n13458), .O(new_n13459));
  nor2 g13266(.a(new_n13459), .b(new_n13457), .O(new_n13460));
  nor2 g13267(.a(new_n13458), .b(new_n13456), .O(new_n13461));
  nor2 g13268(.a(new_n13461), .b(new_n13460), .O(new_n13462));
  inv1 g13269(.a(new_n13462), .O(new_n13463));
  nor2 g13270(.a(new_n13463), .b(new_n13455), .O(new_n13464));
  nor2 g13271(.a(new_n13462), .b(new_n13454), .O(new_n13465));
  nor2 g13272(.a(new_n13465), .b(new_n13464), .O(new_n13466));
  inv1 g13273(.a(new_n13466), .O(new_n13467));
  nor2 g13274(.a(new_n13218), .b(new_n13212), .O(new_n13468));
  nor2 g13275(.a(new_n13010), .b(new_n13003), .O(new_n13469));
  nor2 g13276(.a(new_n13182), .b(new_n13175), .O(new_n13470));
  nor2 g13277(.a(new_n13470), .b(new_n13469), .O(new_n13471));
  inv1 g13278(.a(new_n13469), .O(new_n13472));
  inv1 g13279(.a(new_n13470), .O(new_n13473));
  nor2 g13280(.a(new_n13473), .b(new_n13472), .O(new_n13474));
  nor2 g13281(.a(new_n13474), .b(new_n13471), .O(new_n13475));
  nor2 g13282(.a(new_n13169), .b(new_n13162), .O(new_n13476));
  nor2 g13283(.a(new_n13476), .b(new_n13475), .O(new_n13477));
  inv1 g13284(.a(new_n13475), .O(new_n13478));
  inv1 g13285(.a(new_n13476), .O(new_n13479));
  nor2 g13286(.a(new_n13479), .b(new_n13478), .O(new_n13480));
  nor2 g13287(.a(new_n13480), .b(new_n13477), .O(new_n13481));
  inv1 g13288(.a(new_n13481), .O(new_n13482));
  nor2 g13289(.a(new_n13068), .b(new_n13061), .O(new_n13483));
  nor2 g13290(.a(new_n13123), .b(new_n13116), .O(new_n13484));
  nor2 g13291(.a(new_n13484), .b(new_n13483), .O(new_n13485));
  inv1 g13292(.a(new_n13483), .O(new_n13486));
  inv1 g13293(.a(new_n13484), .O(new_n13487));
  nor2 g13294(.a(new_n13487), .b(new_n13486), .O(new_n13488));
  nor2 g13295(.a(new_n13488), .b(new_n13485), .O(new_n13489));
  nor2 g13296(.a(new_n13157), .b(new_n13151), .O(new_n13490));
  nor2 g13297(.a(new_n13490), .b(new_n13489), .O(new_n13491));
  inv1 g13298(.a(new_n13489), .O(new_n13492));
  inv1 g13299(.a(new_n13490), .O(new_n13493));
  nor2 g13300(.a(new_n13493), .b(new_n13492), .O(new_n13494));
  nor2 g13301(.a(new_n13494), .b(new_n13491), .O(new_n13495));
  inv1 g13302(.a(new_n13495), .O(new_n13496));
  nor2 g13303(.a(new_n13496), .b(new_n13482), .O(new_n13497));
  nor2 g13304(.a(new_n13495), .b(new_n13481), .O(new_n13498));
  nor2 g13305(.a(new_n13498), .b(new_n13497), .O(new_n13499));
  inv1 g13306(.a(new_n13499), .O(new_n13500));
  nor2 g13307(.a(new_n13500), .b(new_n13468), .O(new_n13501));
  inv1 g13308(.a(new_n13468), .O(new_n13502));
  nor2 g13309(.a(new_n13499), .b(new_n13502), .O(new_n13503));
  nor2 g13310(.a(new_n13503), .b(new_n13501), .O(new_n13504));
  inv1 g13311(.a(new_n13504), .O(new_n13505));
  nor2 g13312(.a(new_n13505), .b(new_n13467), .O(new_n13506));
  nor2 g13313(.a(new_n13504), .b(new_n13466), .O(new_n13507));
  nor2 g13314(.a(new_n13507), .b(new_n13506), .O(new_n13508));
  inv1 g13315(.a(new_n13508), .O(new_n13509));
  nor2 g13316(.a(new_n13509), .b(new_n13441), .O(new_n13510));
  inv1 g13317(.a(new_n13441), .O(new_n13511));
  nor2 g13318(.a(new_n13508), .b(new_n13511), .O(new_n13512));
  nor2 g13319(.a(new_n13512), .b(new_n13510), .O(new_n13513));
  inv1 g13320(.a(new_n13513), .O(new_n13514));
  nor2 g13321(.a(new_n12982), .b(new_n12978), .O(new_n13515));
  nor2 g13322(.a(new_n13198), .b(new_n13194), .O(new_n13516));
  nor2 g13323(.a(new_n12953), .b(new_n12947), .O(new_n13517));
  inv1 g13324(.a(new_n13517), .O(new_n13518));
  nor2 g13325(.a(new_n13013), .b(new_n12993), .O(new_n13519));
  nor2 g13326(.a(new_n13519), .b(new_n13518), .O(new_n13520));
  inv1 g13327(.a(new_n13519), .O(new_n13521));
  nor2 g13328(.a(new_n13521), .b(new_n13517), .O(new_n13522));
  nor2 g13329(.a(new_n13522), .b(new_n13520), .O(new_n13523));
  nor2 g13330(.a(new_n13191), .b(new_n13184), .O(new_n13524));
  inv1 g13331(.a(new_n13524), .O(new_n13525));
  nor2 g13332(.a(new_n13525), .b(new_n13523), .O(new_n13526));
  inv1 g13333(.a(new_n13523), .O(new_n13527));
  nor2 g13334(.a(new_n13524), .b(new_n13527), .O(new_n13528));
  nor2 g13335(.a(new_n13528), .b(new_n13526), .O(new_n13529));
  inv1 g13336(.a(new_n13529), .O(new_n13530));
  nor2 g13337(.a(new_n12967), .b(new_n12960), .O(new_n13531));
  inv1 g13338(.a(new_n13531), .O(new_n13532));
  nor2 g13339(.a(new_n10468), .b(new_n322), .O(new_n13533));
  nor2 g13340(.a(new_n10895), .b(new_n295), .O(new_n13534));
  nor2 g13341(.a(new_n13534), .b(new_n13533), .O(new_n13535));
  nor2 g13342(.a(new_n10895), .b(new_n322), .O(new_n13536));
  inv1 g13343(.a(new_n13536), .O(new_n13537));
  nor2 g13344(.a(new_n13537), .b(new_n13170), .O(new_n13538));
  nor2 g13345(.a(new_n13538), .b(new_n13535), .O(new_n13539));
  inv1 g13346(.a(new_n13539), .O(new_n13540));
  nor2 g13347(.a(new_n13540), .b(new_n13133), .O(new_n13541));
  nor2 g13348(.a(new_n13539), .b(new_n13134), .O(new_n13542));
  nor2 g13349(.a(new_n13542), .b(new_n13541), .O(new_n13543));
  nor2 g13350(.a(new_n13543), .b(new_n13532), .O(new_n13544));
  inv1 g13351(.a(new_n13543), .O(new_n13545));
  nor2 g13352(.a(new_n13545), .b(new_n13531), .O(new_n13546));
  nor2 g13353(.a(new_n13546), .b(new_n13544), .O(new_n13547));
  nor2 g13354(.a(new_n12939), .b(new_n12933), .O(new_n13548));
  inv1 g13355(.a(new_n13548), .O(new_n13549));
  nor2 g13356(.a(new_n13549), .b(new_n13547), .O(new_n13550));
  inv1 g13357(.a(new_n13547), .O(new_n13551));
  nor2 g13358(.a(new_n13548), .b(new_n13551), .O(new_n13552));
  nor2 g13359(.a(new_n13552), .b(new_n13550), .O(new_n13553));
  inv1 g13360(.a(new_n13553), .O(new_n13554));
  nor2 g13361(.a(new_n13554), .b(new_n13530), .O(new_n13555));
  nor2 g13362(.a(new_n13553), .b(new_n13529), .O(new_n13556));
  nor2 g13363(.a(new_n13556), .b(new_n13555), .O(new_n13557));
  inv1 g13364(.a(new_n13557), .O(new_n13558));
  nor2 g13365(.a(new_n13558), .b(new_n13516), .O(new_n13559));
  inv1 g13366(.a(new_n13516), .O(new_n13560));
  nor2 g13367(.a(new_n13557), .b(new_n13560), .O(new_n13561));
  nor2 g13368(.a(new_n13561), .b(new_n13559), .O(new_n13562));
  inv1 g13369(.a(new_n13562), .O(new_n13563));
  nor2 g13370(.a(new_n13563), .b(new_n13515), .O(new_n13564));
  inv1 g13371(.a(new_n13515), .O(new_n13565));
  nor2 g13372(.a(new_n13562), .b(new_n13565), .O(new_n13566));
  nor2 g13373(.a(new_n13566), .b(new_n13564), .O(new_n13567));
  inv1 g13374(.a(new_n13567), .O(new_n13568));
  nor2 g13375(.a(new_n13568), .b(new_n13514), .O(new_n13569));
  nor2 g13376(.a(new_n13567), .b(new_n13513), .O(new_n13570));
  nor2 g13377(.a(new_n13570), .b(new_n13569), .O(new_n13571));
  inv1 g13378(.a(new_n13571), .O(new_n13572));
  nor2 g13379(.a(new_n13572), .b(new_n13440), .O(new_n13573));
  inv1 g13380(.a(new_n13440), .O(new_n13574));
  nor2 g13381(.a(new_n13571), .b(new_n13574), .O(new_n13575));
  nor2 g13382(.a(new_n13575), .b(new_n13573), .O(new_n13576));
  inv1 g13383(.a(new_n13576), .O(new_n13577));
  nor2 g13384(.a(new_n13577), .b(new_n13439), .O(new_n13578));
  nor2 g13385(.a(new_n13576), .b(new_n13438), .O(new_n13579));
  nor2 g13386(.a(new_n13579), .b(new_n13578), .O(new_n13580));
  nor2 g13387(.a(new_n13580), .b(new_n13257), .O(new_n13581));
  inv1 g13388(.a(new_n13580), .O(new_n13582));
  nor2 g13389(.a(new_n13582), .b(new_n13256), .O(new_n13583));
  nor2 g13390(.a(new_n13583), .b(new_n13581), .O(new_n13584));
  inv1 g13391(.a(new_n13584), .O(new_n13585));
  nor2 g13392(.a(new_n13251), .b(new_n13247), .O(new_n13586));
  nor2 g13393(.a(new_n13586), .b(new_n13585), .O(new_n13587));
  inv1 g13394(.a(new_n13586), .O(new_n13588));
  nor2 g13395(.a(new_n13588), .b(new_n13584), .O(new_n13589));
  nor2 g13396(.a(new_n13589), .b(new_n13587), .O(new_n13590));
  inv1 g13397(.a(new_n13590), .O(\asquared[69] ));
  nor2 g13398(.a(new_n13578), .b(new_n13573), .O(new_n13592));
  nor2 g13399(.a(new_n13435), .b(new_n13430), .O(new_n13593));
  nor2 g13400(.a(new_n13510), .b(new_n13506), .O(new_n13594));
  inv1 g13401(.a(new_n13594), .O(new_n13595));
  nor2 g13402(.a(new_n13417), .b(new_n13365), .O(new_n13596));
  nor2 g13403(.a(new_n13501), .b(new_n13497), .O(new_n13597));
  nor2 g13404(.a(new_n13312), .b(new_n13307), .O(new_n13598));
  nor2 g13405(.a(new_n13328), .b(new_n13321), .O(new_n13599));
  nor2 g13406(.a(new_n13599), .b(new_n13598), .O(new_n13600));
  inv1 g13407(.a(new_n13598), .O(new_n13601));
  inv1 g13408(.a(new_n13599), .O(new_n13602));
  nor2 g13409(.a(new_n13602), .b(new_n13601), .O(new_n13603));
  nor2 g13410(.a(new_n13603), .b(new_n13600), .O(new_n13604));
  nor2 g13411(.a(new_n13405), .b(new_n13397), .O(new_n13605));
  nor2 g13412(.a(new_n13605), .b(new_n13604), .O(new_n13606));
  inv1 g13413(.a(new_n13604), .O(new_n13607));
  inv1 g13414(.a(new_n13605), .O(new_n13608));
  nor2 g13415(.a(new_n13608), .b(new_n13607), .O(new_n13609));
  nor2 g13416(.a(new_n13609), .b(new_n13606), .O(new_n13610));
  inv1 g13417(.a(new_n13610), .O(new_n13611));
  nor2 g13418(.a(new_n13494), .b(new_n13488), .O(new_n13612));
  inv1 g13419(.a(new_n13612), .O(new_n13613));
  nor2 g13420(.a(new_n13453), .b(new_n13447), .O(new_n13614));
  inv1 g13421(.a(new_n13614), .O(new_n13615));
  nor2 g13422(.a(new_n13615), .b(new_n13613), .O(new_n13616));
  nor2 g13423(.a(new_n13614), .b(new_n13612), .O(new_n13617));
  nor2 g13424(.a(new_n13617), .b(new_n13616), .O(new_n13618));
  inv1 g13425(.a(new_n13618), .O(new_n13619));
  nor2 g13426(.a(new_n13619), .b(new_n13611), .O(new_n13620));
  nor2 g13427(.a(new_n13618), .b(new_n13610), .O(new_n13621));
  nor2 g13428(.a(new_n13621), .b(new_n13620), .O(new_n13622));
  inv1 g13429(.a(new_n13622), .O(new_n13623));
  nor2 g13430(.a(new_n13623), .b(new_n13597), .O(new_n13624));
  inv1 g13431(.a(new_n13597), .O(new_n13625));
  nor2 g13432(.a(new_n13622), .b(new_n13625), .O(new_n13626));
  nor2 g13433(.a(new_n13626), .b(new_n13624), .O(new_n13627));
  inv1 g13434(.a(new_n13627), .O(new_n13628));
  nor2 g13435(.a(new_n13628), .b(new_n13596), .O(new_n13629));
  inv1 g13436(.a(new_n13596), .O(new_n13630));
  nor2 g13437(.a(new_n13627), .b(new_n13630), .O(new_n13631));
  nor2 g13438(.a(new_n13631), .b(new_n13629), .O(new_n13632));
  nor2 g13439(.a(new_n13632), .b(new_n13595), .O(new_n13633));
  inv1 g13440(.a(new_n13632), .O(new_n13634));
  nor2 g13441(.a(new_n13634), .b(new_n13594), .O(new_n13635));
  nor2 g13442(.a(new_n13635), .b(new_n13633), .O(new_n13636));
  inv1 g13443(.a(new_n13636), .O(new_n13637));
  nor2 g13444(.a(new_n13272), .b(new_n13266), .O(new_n13638));
  inv1 g13445(.a(new_n13638), .O(new_n13639));
  nor2 g13446(.a(new_n13314), .b(new_n13299), .O(new_n13640));
  inv1 g13447(.a(new_n13640), .O(new_n13641));
  nor2 g13448(.a(new_n13362), .b(new_n13355), .O(new_n13642));
  inv1 g13449(.a(new_n13642), .O(new_n13643));
  nor2 g13450(.a(new_n13643), .b(new_n13641), .O(new_n13644));
  nor2 g13451(.a(new_n13642), .b(new_n13640), .O(new_n13645));
  nor2 g13452(.a(new_n13645), .b(new_n13644), .O(new_n13646));
  nor2 g13453(.a(new_n13552), .b(new_n13546), .O(new_n13647));
  inv1 g13454(.a(new_n13647), .O(new_n13648));
  nor2 g13455(.a(new_n13648), .b(new_n13646), .O(new_n13649));
  inv1 g13456(.a(new_n13646), .O(new_n13650));
  nor2 g13457(.a(new_n13647), .b(new_n13650), .O(new_n13651));
  nor2 g13458(.a(new_n13651), .b(new_n13649), .O(new_n13652));
  inv1 g13459(.a(new_n13652), .O(new_n13653));
  nor2 g13460(.a(new_n13380), .b(new_n13373), .O(new_n13654));
  nor2 g13461(.a(new_n13391), .b(new_n13385), .O(new_n13655));
  nor2 g13462(.a(new_n13655), .b(new_n13654), .O(new_n13656));
  inv1 g13463(.a(new_n13654), .O(new_n13657));
  inv1 g13464(.a(new_n13655), .O(new_n13658));
  nor2 g13465(.a(new_n13658), .b(new_n13657), .O(new_n13659));
  nor2 g13466(.a(new_n13659), .b(new_n13656), .O(new_n13660));
  nor2 g13467(.a(new_n13353), .b(new_n13346), .O(new_n13661));
  nor2 g13468(.a(new_n13661), .b(new_n13660), .O(new_n13662));
  inv1 g13469(.a(new_n13660), .O(new_n13663));
  inv1 g13470(.a(new_n13661), .O(new_n13664));
  nor2 g13471(.a(new_n13664), .b(new_n13663), .O(new_n13665));
  nor2 g13472(.a(new_n13665), .b(new_n13662), .O(new_n13666));
  inv1 g13473(.a(new_n13666), .O(new_n13667));
  nor2 g13474(.a(new_n13297), .b(new_n13290), .O(new_n13668));
  nor2 g13475(.a(new_n13283), .b(new_n13277), .O(new_n13669));
  nor2 g13476(.a(new_n13669), .b(new_n13668), .O(new_n13670));
  inv1 g13477(.a(new_n13668), .O(new_n13671));
  inv1 g13478(.a(new_n13669), .O(new_n13672));
  nor2 g13479(.a(new_n13672), .b(new_n13671), .O(new_n13673));
  nor2 g13480(.a(new_n13673), .b(new_n13670), .O(new_n13674));
  nor2 g13481(.a(new_n13338), .b(new_n13332), .O(new_n13675));
  nor2 g13482(.a(new_n13675), .b(new_n13674), .O(new_n13676));
  inv1 g13483(.a(new_n13674), .O(new_n13677));
  inv1 g13484(.a(new_n13675), .O(new_n13678));
  nor2 g13485(.a(new_n13678), .b(new_n13677), .O(new_n13679));
  nor2 g13486(.a(new_n13679), .b(new_n13676), .O(new_n13680));
  nor2 g13487(.a(new_n13414), .b(new_n13407), .O(new_n13681));
  inv1 g13488(.a(new_n13681), .O(new_n13682));
  nor2 g13489(.a(new_n13682), .b(new_n13680), .O(new_n13683));
  inv1 g13490(.a(new_n13680), .O(new_n13684));
  nor2 g13491(.a(new_n13681), .b(new_n13684), .O(new_n13685));
  nor2 g13492(.a(new_n13685), .b(new_n13683), .O(new_n13686));
  inv1 g13493(.a(new_n13686), .O(new_n13687));
  nor2 g13494(.a(new_n13687), .b(new_n13667), .O(new_n13688));
  nor2 g13495(.a(new_n13686), .b(new_n13666), .O(new_n13689));
  nor2 g13496(.a(new_n13689), .b(new_n13688), .O(new_n13690));
  inv1 g13497(.a(new_n13690), .O(new_n13691));
  nor2 g13498(.a(new_n13691), .b(new_n13653), .O(new_n13692));
  nor2 g13499(.a(new_n13690), .b(new_n13652), .O(new_n13693));
  nor2 g13500(.a(new_n13693), .b(new_n13692), .O(new_n13694));
  nor2 g13501(.a(new_n13694), .b(new_n13639), .O(new_n13695));
  inv1 g13502(.a(new_n13694), .O(new_n13696));
  nor2 g13503(.a(new_n13696), .b(new_n13638), .O(new_n13697));
  nor2 g13504(.a(new_n13697), .b(new_n13695), .O(new_n13698));
  inv1 g13505(.a(new_n13698), .O(new_n13699));
  nor2 g13506(.a(new_n13699), .b(new_n13637), .O(new_n13700));
  nor2 g13507(.a(new_n13698), .b(new_n13636), .O(new_n13701));
  nor2 g13508(.a(new_n13701), .b(new_n13700), .O(new_n13702));
  inv1 g13509(.a(new_n13702), .O(new_n13703));
  nor2 g13510(.a(new_n13703), .b(new_n13593), .O(new_n13704));
  inv1 g13511(.a(new_n13593), .O(new_n13705));
  nor2 g13512(.a(new_n13702), .b(new_n13705), .O(new_n13706));
  nor2 g13513(.a(new_n13706), .b(new_n13704), .O(new_n13707));
  inv1 g13514(.a(new_n13707), .O(new_n13708));
  nor2 g13515(.a(new_n13569), .b(new_n13564), .O(new_n13709));
  inv1 g13516(.a(new_n13709), .O(new_n13710));
  nor2 g13517(.a(new_n13425), .b(new_n13421), .O(new_n13711));
  inv1 g13518(.a(new_n13711), .O(new_n13712));
  nor2 g13519(.a(new_n13712), .b(new_n13710), .O(new_n13713));
  nor2 g13520(.a(new_n13711), .b(new_n13709), .O(new_n13714));
  nor2 g13521(.a(new_n13714), .b(new_n13713), .O(new_n13715));
  inv1 g13522(.a(new_n13715), .O(new_n13716));
  nor2 g13523(.a(new_n13528), .b(new_n13522), .O(new_n13717));
  inv1 g13524(.a(new_n13717), .O(new_n13718));
  nor2 g13525(.a(new_n5178), .b(new_n2184), .O(new_n13719));
  nor2 g13526(.a(new_n13719), .b(new_n13322), .O(new_n13720));
  inv1 g13527(.a(new_n13320), .O(new_n13721));
  nor2 g13528(.a(new_n5393), .b(new_n2184), .O(new_n13722));
  inv1 g13529(.a(new_n13722), .O(new_n13723));
  nor2 g13530(.a(new_n13723), .b(new_n13721), .O(new_n13724));
  nor2 g13531(.a(new_n13724), .b(new_n13720), .O(new_n13725));
  nor2 g13532(.a(new_n13725), .b(new_n13375), .O(new_n13726));
  inv1 g13533(.a(new_n13725), .O(new_n13727));
  nor2 g13534(.a(new_n13727), .b(new_n13374), .O(new_n13728));
  nor2 g13535(.a(new_n13728), .b(new_n13726), .O(new_n13729));
  inv1 g13536(.a(new_n13729), .O(new_n13730));
  nor2 g13537(.a(new_n10468), .b(new_n363), .O(new_n13731));
  nor2 g13538(.a(new_n10320), .b(new_n438), .O(new_n13732));
  nor2 g13539(.a(new_n13732), .b(new_n13731), .O(new_n13733));
  nor2 g13540(.a(new_n10468), .b(new_n438), .O(new_n13734));
  inv1 g13541(.a(new_n13734), .O(new_n13735));
  nor2 g13542(.a(new_n13735), .b(new_n13165), .O(new_n13736));
  nor2 g13543(.a(new_n13736), .b(new_n13733), .O(new_n13737));
  inv1 g13544(.a(new_n13737), .O(new_n13738));
  nor2 g13545(.a(new_n13738), .b(new_n13536), .O(new_n13739));
  nor2 g13546(.a(new_n13737), .b(new_n13537), .O(new_n13740));
  nor2 g13547(.a(new_n13740), .b(new_n13739), .O(new_n13741));
  nor2 g13548(.a(new_n5971), .b(new_n1736), .O(new_n13742));
  nor2 g13549(.a(new_n5796), .b(new_n1903), .O(new_n13743));
  nor2 g13550(.a(new_n13743), .b(new_n13742), .O(new_n13744));
  nor2 g13551(.a(new_n5971), .b(new_n1903), .O(new_n13745));
  inv1 g13552(.a(new_n13745), .O(new_n13746));
  nor2 g13553(.a(new_n13746), .b(new_n13177), .O(new_n13747));
  nor2 g13554(.a(new_n13747), .b(new_n13744), .O(new_n13748));
  nor2 g13555(.a(new_n13748), .b(new_n13348), .O(new_n13749));
  inv1 g13556(.a(new_n13748), .O(new_n13750));
  nor2 g13557(.a(new_n13750), .b(new_n13347), .O(new_n13751));
  nor2 g13558(.a(new_n13751), .b(new_n13749), .O(new_n13752));
  nor2 g13559(.a(new_n13752), .b(new_n13741), .O(new_n13753));
  inv1 g13560(.a(new_n13741), .O(new_n13754));
  inv1 g13561(.a(new_n13752), .O(new_n13755));
  nor2 g13562(.a(new_n13755), .b(new_n13754), .O(new_n13756));
  nor2 g13563(.a(new_n13756), .b(new_n13753), .O(new_n13757));
  nor2 g13564(.a(new_n13757), .b(new_n13730), .O(new_n13758));
  inv1 g13565(.a(new_n13757), .O(new_n13759));
  nor2 g13566(.a(new_n13759), .b(new_n13729), .O(new_n13760));
  nor2 g13567(.a(new_n13760), .b(new_n13758), .O(new_n13761));
  nor2 g13568(.a(new_n13761), .b(new_n13718), .O(new_n13762));
  inv1 g13569(.a(new_n13761), .O(new_n13763));
  nor2 g13570(.a(new_n13763), .b(new_n13717), .O(new_n13764));
  nor2 g13571(.a(new_n13764), .b(new_n13762), .O(new_n13765));
  inv1 g13572(.a(new_n13765), .O(new_n13766));
  nor2 g13573(.a(new_n8946), .b(new_n699), .O(new_n13767));
  inv1 g13574(.a(new_n13767), .O(new_n13768));
  nor2 g13575(.a(new_n6893), .b(new_n1425), .O(new_n13769));
  nor2 g13576(.a(new_n6570), .b(new_n1493), .O(new_n13770));
  nor2 g13577(.a(new_n13770), .b(new_n13769), .O(new_n13771));
  nor2 g13578(.a(new_n6893), .b(new_n1493), .O(new_n13772));
  inv1 g13579(.a(new_n13772), .O(new_n13773));
  nor2 g13580(.a(new_n13773), .b(new_n13370), .O(new_n13774));
  nor2 g13581(.a(new_n13774), .b(new_n13771), .O(new_n13775));
  nor2 g13582(.a(new_n13775), .b(new_n13768), .O(new_n13776));
  inv1 g13583(.a(new_n13775), .O(new_n13777));
  nor2 g13584(.a(new_n13777), .b(new_n13767), .O(new_n13778));
  nor2 g13585(.a(new_n13778), .b(new_n13776), .O(new_n13779));
  nor2 g13586(.a(new_n9156), .b(new_n613), .O(new_n13780));
  nor2 g13587(.a(new_n9658), .b(new_n569), .O(new_n13781));
  nor2 g13588(.a(new_n13781), .b(new_n13780), .O(new_n13782));
  nor2 g13589(.a(new_n9658), .b(new_n613), .O(new_n13783));
  inv1 g13590(.a(new_n13783), .O(new_n13784));
  nor2 g13591(.a(new_n13784), .b(new_n13306), .O(new_n13785));
  nor2 g13592(.a(new_n13785), .b(new_n13782), .O(new_n13786));
  nor2 g13593(.a(new_n13786), .b(new_n13387), .O(new_n13787));
  inv1 g13594(.a(new_n13786), .O(new_n13788));
  nor2 g13595(.a(new_n13788), .b(new_n13386), .O(new_n13789));
  nor2 g13596(.a(new_n13789), .b(new_n13787), .O(new_n13790));
  nor2 g13597(.a(new_n13541), .b(new_n13538), .O(new_n13791));
  nor2 g13598(.a(new_n13791), .b(new_n13790), .O(new_n13792));
  inv1 g13599(.a(new_n13790), .O(new_n13793));
  inv1 g13600(.a(new_n13791), .O(new_n13794));
  nor2 g13601(.a(new_n13794), .b(new_n13793), .O(new_n13795));
  nor2 g13602(.a(new_n13795), .b(new_n13792), .O(new_n13796));
  inv1 g13603(.a(new_n13796), .O(new_n13797));
  nor2 g13604(.a(new_n13797), .b(new_n13779), .O(new_n13798));
  inv1 g13605(.a(new_n13779), .O(new_n13799));
  nor2 g13606(.a(new_n13796), .b(new_n13799), .O(new_n13800));
  nor2 g13607(.a(new_n13800), .b(new_n13798), .O(new_n13801));
  inv1 g13608(.a(new_n13801), .O(new_n13802));
  nor2 g13609(.a(new_n13802), .b(new_n13766), .O(new_n13803));
  nor2 g13610(.a(new_n13801), .b(new_n13765), .O(new_n13804));
  nor2 g13611(.a(new_n13804), .b(new_n13803), .O(new_n13805));
  inv1 g13612(.a(new_n13805), .O(new_n13806));
  nor2 g13613(.a(new_n13559), .b(new_n13555), .O(new_n13807));
  nor2 g13614(.a(new_n13464), .b(new_n13461), .O(new_n13808));
  nor2 g13615(.a(new_n13480), .b(new_n13474), .O(new_n13809));
  inv1 g13616(.a(new_n13809), .O(new_n13810));
  nor2 g13617(.a(new_n11046), .b(new_n9318), .O(new_n13811));
  nor2 g13618(.a(new_n10280), .b(new_n9506), .O(new_n13812));
  nor2 g13619(.a(new_n13812), .b(new_n13811), .O(new_n13813));
  inv1 g13620(.a(new_n13813), .O(new_n13814));
  nor2 g13621(.a(new_n13814), .b(new_n13278), .O(new_n13815));
  nor2 g13622(.a(new_n13813), .b(new_n13279), .O(new_n13816));
  nor2 g13623(.a(new_n13816), .b(new_n13815), .O(new_n13817));
  nor2 g13624(.a(new_n4954), .b(new_n2433), .O(new_n13818));
  inv1 g13625(.a(new_n13818), .O(new_n13819));
  nor2 g13626(.a(new_n4425), .b(new_n2660), .O(new_n13820));
  nor2 g13627(.a(new_n13820), .b(new_n13399), .O(new_n13821));
  inv1 g13628(.a(new_n13396), .O(new_n13822));
  nor2 g13629(.a(new_n4682), .b(new_n2660), .O(new_n13823));
  inv1 g13630(.a(new_n13823), .O(new_n13824));
  nor2 g13631(.a(new_n13824), .b(new_n13822), .O(new_n13825));
  nor2 g13632(.a(new_n13825), .b(new_n13821), .O(new_n13826));
  nor2 g13633(.a(new_n13826), .b(new_n13819), .O(new_n13827));
  inv1 g13634(.a(new_n13826), .O(new_n13828));
  nor2 g13635(.a(new_n13828), .b(new_n13818), .O(new_n13829));
  nor2 g13636(.a(new_n13829), .b(new_n13827), .O(new_n13830));
  nor2 g13637(.a(new_n13830), .b(new_n13817), .O(new_n13831));
  inv1 g13638(.a(new_n13817), .O(new_n13832));
  inv1 g13639(.a(new_n13830), .O(new_n13833));
  nor2 g13640(.a(new_n13833), .b(new_n13832), .O(new_n13834));
  nor2 g13641(.a(new_n13834), .b(new_n13831), .O(new_n13835));
  nor2 g13642(.a(new_n13835), .b(new_n13810), .O(new_n13836));
  inv1 g13643(.a(new_n13835), .O(new_n13837));
  nor2 g13644(.a(new_n13837), .b(new_n13809), .O(new_n13838));
  nor2 g13645(.a(new_n13838), .b(new_n13836), .O(new_n13839));
  inv1 g13646(.a(new_n13839), .O(new_n13840));
  nor2 g13647(.a(new_n8476), .b(new_n800), .O(new_n13841));
  inv1 g13648(.a(new_n13841), .O(new_n13842));
  nor2 g13649(.a(new_n6958), .b(new_n1297), .O(new_n13843));
  nor2 g13650(.a(new_n13843), .b(new_n13333), .O(new_n13844));
  inv1 g13651(.a(new_n13843), .O(new_n13845));
  nor2 g13652(.a(new_n13845), .b(new_n13334), .O(new_n13846));
  nor2 g13653(.a(new_n13846), .b(new_n13844), .O(new_n13847));
  nor2 g13654(.a(new_n13847), .b(new_n13842), .O(new_n13848));
  inv1 g13655(.a(new_n13847), .O(new_n13849));
  nor2 g13656(.a(new_n13849), .b(new_n13841), .O(new_n13850));
  nor2 g13657(.a(new_n13850), .b(new_n13848), .O(new_n13851));
  inv1 g13658(.a(new_n13851), .O(new_n13852));
  nor2 g13659(.a(new_n4366), .b(new_n2826), .O(new_n13853));
  inv1 g13660(.a(new_n13853), .O(new_n13854));
  nor2 g13661(.a(new_n3870), .b(new_n3231), .O(new_n13855));
  nor2 g13662(.a(new_n13855), .b(new_n13291), .O(new_n13856));
  inv1 g13663(.a(new_n13288), .O(new_n13857));
  nor2 g13664(.a(new_n4093), .b(new_n3231), .O(new_n13858));
  inv1 g13665(.a(new_n13858), .O(new_n13859));
  nor2 g13666(.a(new_n13859), .b(new_n13857), .O(new_n13860));
  nor2 g13667(.a(new_n13860), .b(new_n13856), .O(new_n13861));
  nor2 g13668(.a(new_n13861), .b(new_n13854), .O(new_n13862));
  inv1 g13669(.a(new_n13861), .O(new_n13863));
  nor2 g13670(.a(new_n13863), .b(new_n13853), .O(new_n13864));
  nor2 g13671(.a(new_n13864), .b(new_n13862), .O(new_n13865));
  nor2 g13672(.a(new_n11186), .b(new_n295), .O(new_n13866));
  inv1 g13673(.a(new_n13866), .O(new_n13867));
  nor2 g13674(.a(new_n3722), .b(\a[34] ), .O(new_n13868));
  nor2 g13675(.a(new_n13868), .b(new_n13867), .O(new_n13869));
  inv1 g13676(.a(new_n13868), .O(new_n13870));
  nor2 g13677(.a(new_n13870), .b(new_n13866), .O(new_n13871));
  nor2 g13678(.a(new_n13871), .b(new_n13869), .O(new_n13872));
  nor2 g13679(.a(new_n13872), .b(new_n13865), .O(new_n13873));
  inv1 g13680(.a(new_n13865), .O(new_n13874));
  inv1 g13681(.a(new_n13872), .O(new_n13875));
  nor2 g13682(.a(new_n13875), .b(new_n13874), .O(new_n13876));
  nor2 g13683(.a(new_n13876), .b(new_n13873), .O(new_n13877));
  nor2 g13684(.a(new_n13877), .b(new_n13852), .O(new_n13878));
  inv1 g13685(.a(new_n13877), .O(new_n13879));
  nor2 g13686(.a(new_n13879), .b(new_n13851), .O(new_n13880));
  nor2 g13687(.a(new_n13880), .b(new_n13878), .O(new_n13881));
  inv1 g13688(.a(new_n13881), .O(new_n13882));
  nor2 g13689(.a(new_n13882), .b(new_n13840), .O(new_n13883));
  nor2 g13690(.a(new_n13881), .b(new_n13839), .O(new_n13884));
  nor2 g13691(.a(new_n13884), .b(new_n13883), .O(new_n13885));
  inv1 g13692(.a(new_n13885), .O(new_n13886));
  nor2 g13693(.a(new_n13886), .b(new_n13808), .O(new_n13887));
  inv1 g13694(.a(new_n13808), .O(new_n13888));
  nor2 g13695(.a(new_n13885), .b(new_n13888), .O(new_n13889));
  nor2 g13696(.a(new_n13889), .b(new_n13887), .O(new_n13890));
  inv1 g13697(.a(new_n13890), .O(new_n13891));
  nor2 g13698(.a(new_n13891), .b(new_n13807), .O(new_n13892));
  inv1 g13699(.a(new_n13807), .O(new_n13893));
  nor2 g13700(.a(new_n13890), .b(new_n13893), .O(new_n13894));
  nor2 g13701(.a(new_n13894), .b(new_n13892), .O(new_n13895));
  inv1 g13702(.a(new_n13895), .O(new_n13896));
  nor2 g13703(.a(new_n13896), .b(new_n13806), .O(new_n13897));
  nor2 g13704(.a(new_n13895), .b(new_n13805), .O(new_n13898));
  nor2 g13705(.a(new_n13898), .b(new_n13897), .O(new_n13899));
  inv1 g13706(.a(new_n13899), .O(new_n13900));
  nor2 g13707(.a(new_n13900), .b(new_n13716), .O(new_n13901));
  nor2 g13708(.a(new_n13899), .b(new_n13715), .O(new_n13902));
  nor2 g13709(.a(new_n13902), .b(new_n13901), .O(new_n13903));
  inv1 g13710(.a(new_n13903), .O(new_n13904));
  nor2 g13711(.a(new_n13904), .b(new_n13708), .O(new_n13905));
  nor2 g13712(.a(new_n13903), .b(new_n13707), .O(new_n13906));
  nor2 g13713(.a(new_n13906), .b(new_n13905), .O(new_n13907));
  inv1 g13714(.a(new_n13907), .O(new_n13908));
  nor2 g13715(.a(new_n13908), .b(new_n13592), .O(new_n13909));
  inv1 g13716(.a(new_n13592), .O(new_n13910));
  nor2 g13717(.a(new_n13907), .b(new_n13910), .O(new_n13911));
  nor2 g13718(.a(new_n13911), .b(new_n13909), .O(new_n13912));
  inv1 g13719(.a(new_n13912), .O(new_n13913));
  nor2 g13720(.a(new_n13587), .b(new_n13581), .O(new_n13914));
  nor2 g13721(.a(new_n13914), .b(new_n13913), .O(new_n13915));
  inv1 g13722(.a(new_n13914), .O(new_n13916));
  nor2 g13723(.a(new_n13916), .b(new_n13912), .O(new_n13917));
  nor2 g13724(.a(new_n13917), .b(new_n13915), .O(new_n13918));
  inv1 g13725(.a(new_n13918), .O(\asquared[70] ));
  nor2 g13726(.a(new_n13905), .b(new_n13704), .O(new_n13920));
  inv1 g13727(.a(new_n13920), .O(new_n13921));
  nor2 g13728(.a(new_n13700), .b(new_n13635), .O(new_n13922));
  nor2 g13729(.a(new_n13838), .b(new_n13831), .O(new_n13923));
  inv1 g13730(.a(new_n13923), .O(new_n13924));
  nor2 g13731(.a(new_n13728), .b(new_n13720), .O(new_n13925));
  nor2 g13732(.a(new_n13829), .b(new_n13821), .O(new_n13926));
  nor2 g13733(.a(new_n13926), .b(new_n13925), .O(new_n13927));
  inv1 g13734(.a(new_n13925), .O(new_n13928));
  inv1 g13735(.a(new_n13926), .O(new_n13929));
  nor2 g13736(.a(new_n13929), .b(new_n13928), .O(new_n13930));
  nor2 g13737(.a(new_n13930), .b(new_n13927), .O(new_n13931));
  nor2 g13738(.a(new_n13751), .b(new_n13744), .O(new_n13932));
  nor2 g13739(.a(new_n13932), .b(new_n13931), .O(new_n13933));
  inv1 g13740(.a(new_n13931), .O(new_n13934));
  inv1 g13741(.a(new_n13932), .O(new_n13935));
  nor2 g13742(.a(new_n13935), .b(new_n13934), .O(new_n13936));
  nor2 g13743(.a(new_n13936), .b(new_n13933), .O(new_n13937));
  inv1 g13744(.a(new_n13937), .O(new_n13938));
  nor2 g13745(.a(new_n11186), .b(new_n322), .O(new_n13939));
  inv1 g13746(.a(new_n13939), .O(new_n13940));
  nor2 g13747(.a(new_n13871), .b(new_n3722), .O(new_n13941));
  inv1 g13748(.a(new_n13941), .O(new_n13942));
  nor2 g13749(.a(new_n13942), .b(new_n13940), .O(new_n13943));
  nor2 g13750(.a(new_n13941), .b(new_n13939), .O(new_n13944));
  nor2 g13751(.a(new_n13944), .b(new_n13943), .O(new_n13945));
  inv1 g13752(.a(new_n13945), .O(new_n13946));
  nor2 g13753(.a(new_n13864), .b(new_n13856), .O(new_n13947));
  inv1 g13754(.a(new_n13947), .O(new_n13948));
  nor2 g13755(.a(new_n13948), .b(new_n13946), .O(new_n13949));
  nor2 g13756(.a(new_n13947), .b(new_n13945), .O(new_n13950));
  nor2 g13757(.a(new_n13950), .b(new_n13949), .O(new_n13951));
  inv1 g13758(.a(new_n13951), .O(new_n13952));
  nor2 g13759(.a(new_n13952), .b(new_n13938), .O(new_n13953));
  nor2 g13760(.a(new_n13951), .b(new_n13937), .O(new_n13954));
  nor2 g13761(.a(new_n13954), .b(new_n13953), .O(new_n13955));
  nor2 g13762(.a(new_n13955), .b(new_n13924), .O(new_n13956));
  inv1 g13763(.a(new_n13955), .O(new_n13957));
  nor2 g13764(.a(new_n13957), .b(new_n13923), .O(new_n13958));
  nor2 g13765(.a(new_n13958), .b(new_n13956), .O(new_n13959));
  nor2 g13766(.a(new_n13887), .b(new_n13883), .O(new_n13960));
  nor2 g13767(.a(new_n13798), .b(new_n13792), .O(new_n13961));
  inv1 g13768(.a(new_n13961), .O(new_n13962));
  nor2 g13769(.a(new_n13760), .b(new_n13753), .O(new_n13963));
  inv1 g13770(.a(new_n13963), .O(new_n13964));
  nor2 g13771(.a(new_n13964), .b(new_n13962), .O(new_n13965));
  nor2 g13772(.a(new_n13963), .b(new_n13961), .O(new_n13966));
  nor2 g13773(.a(new_n13966), .b(new_n13965), .O(new_n13967));
  nor2 g13774(.a(new_n13880), .b(new_n13873), .O(new_n13968));
  inv1 g13775(.a(new_n13968), .O(new_n13969));
  nor2 g13776(.a(new_n13969), .b(new_n13967), .O(new_n13970));
  inv1 g13777(.a(new_n13967), .O(new_n13971));
  nor2 g13778(.a(new_n13968), .b(new_n13971), .O(new_n13972));
  nor2 g13779(.a(new_n13972), .b(new_n13970), .O(new_n13973));
  inv1 g13780(.a(new_n13973), .O(new_n13974));
  nor2 g13781(.a(new_n13974), .b(new_n13960), .O(new_n13975));
  inv1 g13782(.a(new_n13960), .O(new_n13976));
  nor2 g13783(.a(new_n13973), .b(new_n13976), .O(new_n13977));
  nor2 g13784(.a(new_n13977), .b(new_n13975), .O(new_n13978));
  nor2 g13785(.a(new_n13978), .b(new_n13959), .O(new_n13979));
  inv1 g13786(.a(new_n13959), .O(new_n13980));
  inv1 g13787(.a(new_n13978), .O(new_n13981));
  nor2 g13788(.a(new_n13981), .b(new_n13980), .O(new_n13982));
  nor2 g13789(.a(new_n13982), .b(new_n13979), .O(new_n13983));
  inv1 g13790(.a(new_n13983), .O(new_n13984));
  nor2 g13791(.a(new_n13984), .b(new_n13922), .O(new_n13985));
  inv1 g13792(.a(new_n13922), .O(new_n13986));
  nor2 g13793(.a(new_n13983), .b(new_n13986), .O(new_n13987));
  nor2 g13794(.a(new_n13987), .b(new_n13985), .O(new_n13988));
  inv1 g13795(.a(new_n13988), .O(new_n13989));
  nor2 g13796(.a(new_n13629), .b(new_n13624), .O(new_n13990));
  nor2 g13797(.a(new_n13620), .b(new_n13617), .O(new_n13991));
  nor2 g13798(.a(new_n13850), .b(new_n13844), .O(new_n13992));
  nor2 g13799(.a(new_n13815), .b(new_n13811), .O(new_n13993));
  nor2 g13800(.a(new_n13993), .b(new_n13992), .O(new_n13994));
  inv1 g13801(.a(new_n13992), .O(new_n13995));
  inv1 g13802(.a(new_n13993), .O(new_n13996));
  nor2 g13803(.a(new_n13996), .b(new_n13995), .O(new_n13997));
  nor2 g13804(.a(new_n13997), .b(new_n13994), .O(new_n13998));
  inv1 g13805(.a(new_n13998), .O(new_n13999));
  nor2 g13806(.a(new_n4366), .b(new_n3057), .O(new_n14000));
  inv1 g13807(.a(new_n14000), .O(new_n14001));
  nor2 g13808(.a(new_n3870), .b(new_n3533), .O(new_n14002));
  nor2 g13809(.a(new_n14002), .b(new_n13858), .O(new_n14003));
  inv1 g13810(.a(new_n13855), .O(new_n14004));
  nor2 g13811(.a(new_n4093), .b(new_n3533), .O(new_n14005));
  inv1 g13812(.a(new_n14005), .O(new_n14006));
  nor2 g13813(.a(new_n14006), .b(new_n14004), .O(new_n14007));
  nor2 g13814(.a(new_n14007), .b(new_n14003), .O(new_n14008));
  nor2 g13815(.a(new_n14008), .b(new_n14001), .O(new_n14009));
  inv1 g13816(.a(new_n14008), .O(new_n14010));
  nor2 g13817(.a(new_n14010), .b(new_n14000), .O(new_n14011));
  nor2 g13818(.a(new_n14011), .b(new_n14009), .O(new_n14012));
  inv1 g13819(.a(new_n14012), .O(new_n14013));
  nor2 g13820(.a(new_n14013), .b(new_n13999), .O(new_n14014));
  nor2 g13821(.a(new_n14012), .b(new_n13998), .O(new_n14015));
  nor2 g13822(.a(new_n14015), .b(new_n14014), .O(new_n14016));
  nor2 g13823(.a(new_n14016), .b(new_n13991), .O(new_n14017));
  inv1 g13824(.a(new_n13991), .O(new_n14018));
  inv1 g13825(.a(new_n14016), .O(new_n14019));
  nor2 g13826(.a(new_n14019), .b(new_n14018), .O(new_n14020));
  nor2 g13827(.a(new_n14020), .b(new_n14017), .O(new_n14021));
  inv1 g13828(.a(new_n14021), .O(new_n14022));
  nor2 g13829(.a(new_n9873), .b(new_n569), .O(new_n14023));
  inv1 g13830(.a(new_n14023), .O(new_n14024));
  nor2 g13831(.a(new_n13783), .b(new_n6619), .O(new_n14025));
  nor2 g13832(.a(new_n12580), .b(new_n9518), .O(new_n14026));
  nor2 g13833(.a(new_n14026), .b(new_n14025), .O(new_n14027));
  nor2 g13834(.a(new_n14027), .b(new_n14024), .O(new_n14028));
  inv1 g13835(.a(new_n14027), .O(new_n14029));
  nor2 g13836(.a(new_n14029), .b(new_n14023), .O(new_n14030));
  nor2 g13837(.a(new_n14030), .b(new_n14028), .O(new_n14031));
  inv1 g13838(.a(new_n14031), .O(new_n14032));
  nor2 g13839(.a(new_n10895), .b(new_n363), .O(new_n14033));
  nor2 g13840(.a(new_n10320), .b(new_n502), .O(new_n14034));
  nor2 g13841(.a(new_n14034), .b(new_n13734), .O(new_n14035));
  inv1 g13842(.a(new_n13732), .O(new_n14036));
  nor2 g13843(.a(new_n10468), .b(new_n502), .O(new_n14037));
  inv1 g13844(.a(new_n14037), .O(new_n14038));
  nor2 g13845(.a(new_n14038), .b(new_n14036), .O(new_n14039));
  nor2 g13846(.a(new_n14039), .b(new_n14035), .O(new_n14040));
  inv1 g13847(.a(new_n14040), .O(new_n14041));
  nor2 g13848(.a(new_n14041), .b(new_n14033), .O(new_n14042));
  inv1 g13849(.a(new_n14033), .O(new_n14043));
  nor2 g13850(.a(new_n14040), .b(new_n14043), .O(new_n14044));
  nor2 g13851(.a(new_n14044), .b(new_n14042), .O(new_n14045));
  nor2 g13852(.a(new_n8170), .b(new_n941), .O(new_n14046));
  nor2 g13853(.a(new_n8476), .b(new_n847), .O(new_n14047));
  nor2 g13854(.a(new_n14047), .b(new_n14046), .O(new_n14048));
  nor2 g13855(.a(new_n13334), .b(new_n11665), .O(new_n14049));
  nor2 g13856(.a(new_n14049), .b(new_n14048), .O(new_n14050));
  nor2 g13857(.a(new_n14050), .b(new_n10280), .O(new_n14051));
  inv1 g13858(.a(new_n14050), .O(new_n14052));
  nor2 g13859(.a(new_n14052), .b(new_n10279), .O(new_n14053));
  nor2 g13860(.a(new_n14053), .b(new_n14051), .O(new_n14054));
  nor2 g13861(.a(new_n14054), .b(new_n14045), .O(new_n14055));
  inv1 g13862(.a(new_n14045), .O(new_n14056));
  inv1 g13863(.a(new_n14054), .O(new_n14057));
  nor2 g13864(.a(new_n14057), .b(new_n14056), .O(new_n14058));
  nor2 g13865(.a(new_n14058), .b(new_n14055), .O(new_n14059));
  nor2 g13866(.a(new_n14059), .b(new_n14032), .O(new_n14060));
  inv1 g13867(.a(new_n14059), .O(new_n14061));
  nor2 g13868(.a(new_n14061), .b(new_n14031), .O(new_n14062));
  nor2 g13869(.a(new_n14062), .b(new_n14060), .O(new_n14063));
  inv1 g13870(.a(new_n14063), .O(new_n14064));
  nor2 g13871(.a(new_n14064), .b(new_n14022), .O(new_n14065));
  nor2 g13872(.a(new_n14063), .b(new_n14021), .O(new_n14066));
  nor2 g13873(.a(new_n14066), .b(new_n14065), .O(new_n14067));
  inv1 g13874(.a(new_n14067), .O(new_n14068));
  nor2 g13875(.a(new_n14068), .b(new_n13990), .O(new_n14069));
  inv1 g13876(.a(new_n13990), .O(new_n14070));
  nor2 g13877(.a(new_n14067), .b(new_n14070), .O(new_n14071));
  nor2 g13878(.a(new_n14071), .b(new_n14069), .O(new_n14072));
  inv1 g13879(.a(new_n14072), .O(new_n14073));
  nor2 g13880(.a(new_n13688), .b(new_n13685), .O(new_n14074));
  nor2 g13881(.a(new_n13679), .b(new_n13673), .O(new_n14075));
  inv1 g13882(.a(new_n14075), .O(new_n14076));
  nor2 g13883(.a(new_n4954), .b(new_n2506), .O(new_n14077));
  inv1 g13884(.a(new_n14077), .O(new_n14078));
  nor2 g13885(.a(new_n4425), .b(new_n2826), .O(new_n14079));
  nor2 g13886(.a(new_n14079), .b(new_n13823), .O(new_n14080));
  inv1 g13887(.a(new_n13820), .O(new_n14081));
  nor2 g13888(.a(new_n4682), .b(new_n2826), .O(new_n14082));
  inv1 g13889(.a(new_n14082), .O(new_n14083));
  nor2 g13890(.a(new_n14083), .b(new_n14081), .O(new_n14084));
  nor2 g13891(.a(new_n14084), .b(new_n14080), .O(new_n14085));
  nor2 g13892(.a(new_n14085), .b(new_n14078), .O(new_n14086));
  inv1 g13893(.a(new_n14085), .O(new_n14087));
  nor2 g13894(.a(new_n14087), .b(new_n14077), .O(new_n14088));
  nor2 g13895(.a(new_n14088), .b(new_n14086), .O(new_n14089));
  nor2 g13896(.a(new_n5178), .b(new_n2433), .O(new_n14090));
  inv1 g13897(.a(new_n14090), .O(new_n14091));
  nor2 g13898(.a(new_n6570), .b(new_n1647), .O(new_n14092));
  nor2 g13899(.a(new_n11596), .b(new_n295), .O(new_n14093));
  nor2 g13900(.a(new_n14093), .b(new_n14092), .O(new_n14094));
  inv1 g13901(.a(new_n14092), .O(new_n14095));
  inv1 g13902(.a(new_n14093), .O(new_n14096));
  nor2 g13903(.a(new_n14096), .b(new_n14095), .O(new_n14097));
  nor2 g13904(.a(new_n14097), .b(new_n14094), .O(new_n14098));
  inv1 g13905(.a(new_n14098), .O(new_n14099));
  nor2 g13906(.a(new_n14099), .b(new_n14091), .O(new_n14100));
  nor2 g13907(.a(new_n14098), .b(new_n14090), .O(new_n14101));
  nor2 g13908(.a(new_n14101), .b(new_n14100), .O(new_n14102));
  inv1 g13909(.a(new_n14102), .O(new_n14103));
  nor2 g13910(.a(new_n14103), .b(new_n14089), .O(new_n14104));
  inv1 g13911(.a(new_n14089), .O(new_n14105));
  nor2 g13912(.a(new_n14102), .b(new_n14105), .O(new_n14106));
  nor2 g13913(.a(new_n14106), .b(new_n14104), .O(new_n14107));
  nor2 g13914(.a(new_n14107), .b(new_n14076), .O(new_n14108));
  inv1 g13915(.a(new_n14107), .O(new_n14109));
  nor2 g13916(.a(new_n14109), .b(new_n14075), .O(new_n14110));
  nor2 g13917(.a(new_n14110), .b(new_n14108), .O(new_n14111));
  inv1 g13918(.a(new_n14111), .O(new_n14112));
  nor2 g13919(.a(new_n6958), .b(new_n1425), .O(new_n14113));
  inv1 g13920(.a(new_n14113), .O(new_n14114));
  nor2 g13921(.a(new_n7537), .b(new_n1199), .O(new_n14115));
  nor2 g13922(.a(new_n7294), .b(new_n1297), .O(new_n14116));
  nor2 g13923(.a(new_n14116), .b(new_n14115), .O(new_n14117));
  nor2 g13924(.a(new_n7537), .b(new_n1297), .O(new_n14118));
  inv1 g13925(.a(new_n14118), .O(new_n14119));
  nor2 g13926(.a(new_n14119), .b(new_n13279), .O(new_n14120));
  nor2 g13927(.a(new_n14120), .b(new_n14117), .O(new_n14121));
  nor2 g13928(.a(new_n14121), .b(new_n14114), .O(new_n14122));
  inv1 g13929(.a(new_n14121), .O(new_n14123));
  nor2 g13930(.a(new_n14123), .b(new_n14113), .O(new_n14124));
  nor2 g13931(.a(new_n14124), .b(new_n14122), .O(new_n14125));
  inv1 g13932(.a(new_n14125), .O(new_n14126));
  nor2 g13933(.a(new_n9156), .b(new_n699), .O(new_n14127));
  nor2 g13934(.a(new_n8946), .b(new_n800), .O(new_n14128));
  nor2 g13935(.a(new_n14128), .b(new_n14127), .O(new_n14129));
  nor2 g13936(.a(new_n9156), .b(new_n800), .O(new_n14130));
  inv1 g13937(.a(new_n14130), .O(new_n14131));
  nor2 g13938(.a(new_n14131), .b(new_n13768), .O(new_n14132));
  nor2 g13939(.a(new_n14132), .b(new_n14129), .O(new_n14133));
  inv1 g13940(.a(new_n14133), .O(new_n14134));
  nor2 g13941(.a(new_n14134), .b(new_n13772), .O(new_n14135));
  nor2 g13942(.a(new_n14133), .b(new_n13773), .O(new_n14136));
  nor2 g13943(.a(new_n14136), .b(new_n14135), .O(new_n14137));
  nor2 g13944(.a(new_n5796), .b(new_n2121), .O(new_n14138));
  nor2 g13945(.a(new_n14138), .b(new_n13722), .O(new_n14139));
  nor2 g13946(.a(new_n5796), .b(new_n2184), .O(new_n14140));
  inv1 g13947(.a(new_n14140), .O(new_n14141));
  nor2 g13948(.a(new_n14141), .b(new_n13323), .O(new_n14142));
  nor2 g13949(.a(new_n14142), .b(new_n14139), .O(new_n14143));
  nor2 g13950(.a(new_n14143), .b(new_n13746), .O(new_n14144));
  inv1 g13951(.a(new_n14143), .O(new_n14145));
  nor2 g13952(.a(new_n14145), .b(new_n13745), .O(new_n14146));
  nor2 g13953(.a(new_n14146), .b(new_n14144), .O(new_n14147));
  nor2 g13954(.a(new_n14147), .b(new_n14137), .O(new_n14148));
  inv1 g13955(.a(new_n14137), .O(new_n14149));
  inv1 g13956(.a(new_n14147), .O(new_n14150));
  nor2 g13957(.a(new_n14150), .b(new_n14149), .O(new_n14151));
  nor2 g13958(.a(new_n14151), .b(new_n14148), .O(new_n14152));
  nor2 g13959(.a(new_n14152), .b(new_n14126), .O(new_n14153));
  inv1 g13960(.a(new_n14152), .O(new_n14154));
  nor2 g13961(.a(new_n14154), .b(new_n14125), .O(new_n14155));
  nor2 g13962(.a(new_n14155), .b(new_n14153), .O(new_n14156));
  inv1 g13963(.a(new_n14156), .O(new_n14157));
  nor2 g13964(.a(new_n14157), .b(new_n14112), .O(new_n14158));
  nor2 g13965(.a(new_n14156), .b(new_n14111), .O(new_n14159));
  nor2 g13966(.a(new_n14159), .b(new_n14158), .O(new_n14160));
  inv1 g13967(.a(new_n14160), .O(new_n14161));
  nor2 g13968(.a(new_n14161), .b(new_n14074), .O(new_n14162));
  inv1 g13969(.a(new_n14074), .O(new_n14163));
  nor2 g13970(.a(new_n14160), .b(new_n14163), .O(new_n14164));
  nor2 g13971(.a(new_n14164), .b(new_n14162), .O(new_n14165));
  inv1 g13972(.a(new_n14165), .O(new_n14166));
  nor2 g13973(.a(new_n14166), .b(new_n14073), .O(new_n14167));
  nor2 g13974(.a(new_n14165), .b(new_n14072), .O(new_n14168));
  nor2 g13975(.a(new_n14168), .b(new_n14167), .O(new_n14169));
  inv1 g13976(.a(new_n14169), .O(new_n14170));
  nor2 g13977(.a(new_n14170), .b(new_n13989), .O(new_n14171));
  nor2 g13978(.a(new_n14169), .b(new_n13988), .O(new_n14172));
  nor2 g13979(.a(new_n14172), .b(new_n14171), .O(new_n14173));
  inv1 g13980(.a(new_n14173), .O(new_n14174));
  nor2 g13981(.a(new_n13897), .b(new_n13892), .O(new_n14175));
  inv1 g13982(.a(new_n14175), .O(new_n14176));
  nor2 g13983(.a(new_n13697), .b(new_n13692), .O(new_n14177));
  nor2 g13984(.a(new_n13803), .b(new_n13764), .O(new_n14178));
  nor2 g13985(.a(new_n13651), .b(new_n13645), .O(new_n14179));
  nor2 g13986(.a(new_n13789), .b(new_n13782), .O(new_n14180));
  nor2 g13987(.a(new_n13739), .b(new_n13733), .O(new_n14181));
  nor2 g13988(.a(new_n14181), .b(new_n14180), .O(new_n14182));
  inv1 g13989(.a(new_n14180), .O(new_n14183));
  inv1 g13990(.a(new_n14181), .O(new_n14184));
  nor2 g13991(.a(new_n14184), .b(new_n14183), .O(new_n14185));
  nor2 g13992(.a(new_n14185), .b(new_n14182), .O(new_n14186));
  nor2 g13993(.a(new_n13778), .b(new_n13771), .O(new_n14187));
  nor2 g13994(.a(new_n14187), .b(new_n14186), .O(new_n14188));
  inv1 g13995(.a(new_n14186), .O(new_n14189));
  inv1 g13996(.a(new_n14187), .O(new_n14190));
  nor2 g13997(.a(new_n14190), .b(new_n14189), .O(new_n14191));
  nor2 g13998(.a(new_n14191), .b(new_n14188), .O(new_n14192));
  inv1 g13999(.a(new_n14192), .O(new_n14193));
  nor2 g14000(.a(new_n13665), .b(new_n13659), .O(new_n14194));
  inv1 g14001(.a(new_n14194), .O(new_n14195));
  nor2 g14002(.a(new_n13609), .b(new_n13603), .O(new_n14196));
  inv1 g14003(.a(new_n14196), .O(new_n14197));
  nor2 g14004(.a(new_n14197), .b(new_n14195), .O(new_n14198));
  nor2 g14005(.a(new_n14196), .b(new_n14194), .O(new_n14199));
  nor2 g14006(.a(new_n14199), .b(new_n14198), .O(new_n14200));
  inv1 g14007(.a(new_n14200), .O(new_n14201));
  nor2 g14008(.a(new_n14201), .b(new_n14193), .O(new_n14202));
  nor2 g14009(.a(new_n14200), .b(new_n14192), .O(new_n14203));
  nor2 g14010(.a(new_n14203), .b(new_n14202), .O(new_n14204));
  inv1 g14011(.a(new_n14204), .O(new_n14205));
  nor2 g14012(.a(new_n14205), .b(new_n14179), .O(new_n14206));
  inv1 g14013(.a(new_n14179), .O(new_n14207));
  nor2 g14014(.a(new_n14204), .b(new_n14207), .O(new_n14208));
  nor2 g14015(.a(new_n14208), .b(new_n14206), .O(new_n14209));
  inv1 g14016(.a(new_n14209), .O(new_n14210));
  nor2 g14017(.a(new_n14210), .b(new_n14178), .O(new_n14211));
  inv1 g14018(.a(new_n14178), .O(new_n14212));
  nor2 g14019(.a(new_n14209), .b(new_n14212), .O(new_n14213));
  nor2 g14020(.a(new_n14213), .b(new_n14211), .O(new_n14214));
  inv1 g14021(.a(new_n14214), .O(new_n14215));
  nor2 g14022(.a(new_n14215), .b(new_n14177), .O(new_n14216));
  inv1 g14023(.a(new_n14177), .O(new_n14217));
  nor2 g14024(.a(new_n14214), .b(new_n14217), .O(new_n14218));
  nor2 g14025(.a(new_n14218), .b(new_n14216), .O(new_n14219));
  nor2 g14026(.a(new_n14219), .b(new_n14176), .O(new_n14220));
  inv1 g14027(.a(new_n14219), .O(new_n14221));
  nor2 g14028(.a(new_n14221), .b(new_n14175), .O(new_n14222));
  nor2 g14029(.a(new_n14222), .b(new_n14220), .O(new_n14223));
  inv1 g14030(.a(new_n14223), .O(new_n14224));
  nor2 g14031(.a(new_n13901), .b(new_n13714), .O(new_n14225));
  nor2 g14032(.a(new_n14225), .b(new_n14224), .O(new_n14226));
  inv1 g14033(.a(new_n14225), .O(new_n14227));
  nor2 g14034(.a(new_n14227), .b(new_n14223), .O(new_n14228));
  nor2 g14035(.a(new_n14228), .b(new_n14226), .O(new_n14229));
  inv1 g14036(.a(new_n14229), .O(new_n14230));
  nor2 g14037(.a(new_n14230), .b(new_n14174), .O(new_n14231));
  nor2 g14038(.a(new_n14229), .b(new_n14173), .O(new_n14232));
  nor2 g14039(.a(new_n14232), .b(new_n14231), .O(new_n14233));
  nor2 g14040(.a(new_n14233), .b(new_n13921), .O(new_n14234));
  inv1 g14041(.a(new_n14233), .O(new_n14235));
  nor2 g14042(.a(new_n14235), .b(new_n13920), .O(new_n14236));
  nor2 g14043(.a(new_n14236), .b(new_n14234), .O(new_n14237));
  inv1 g14044(.a(new_n14237), .O(new_n14238));
  nor2 g14045(.a(new_n13915), .b(new_n13911), .O(new_n14239));
  nor2 g14046(.a(new_n14239), .b(new_n14238), .O(new_n14240));
  inv1 g14047(.a(new_n14239), .O(new_n14241));
  nor2 g14048(.a(new_n14241), .b(new_n14237), .O(new_n14242));
  nor2 g14049(.a(new_n14242), .b(new_n14240), .O(new_n14243));
  inv1 g14050(.a(new_n14243), .O(\asquared[71] ));
  nor2 g14051(.a(new_n14231), .b(new_n14226), .O(new_n14245));
  inv1 g14052(.a(new_n14245), .O(new_n14246));
  nor2 g14053(.a(new_n14167), .b(new_n14069), .O(new_n14247));
  inv1 g14054(.a(new_n14247), .O(new_n14248));
  nor2 g14055(.a(new_n13949), .b(new_n13943), .O(new_n14249));
  inv1 g14056(.a(new_n14249), .O(new_n14250));
  nor2 g14057(.a(new_n14014), .b(new_n13994), .O(new_n14251));
  nor2 g14058(.a(new_n14251), .b(new_n14250), .O(new_n14252));
  inv1 g14059(.a(new_n14251), .O(new_n14253));
  nor2 g14060(.a(new_n14253), .b(new_n14249), .O(new_n14254));
  nor2 g14061(.a(new_n14254), .b(new_n14252), .O(new_n14255));
  nor2 g14062(.a(new_n13936), .b(new_n13930), .O(new_n14256));
  inv1 g14063(.a(new_n14256), .O(new_n14257));
  nor2 g14064(.a(new_n14257), .b(new_n14255), .O(new_n14258));
  inv1 g14065(.a(new_n14255), .O(new_n14259));
  nor2 g14066(.a(new_n14256), .b(new_n14259), .O(new_n14260));
  nor2 g14067(.a(new_n14260), .b(new_n14258), .O(new_n14261));
  nor2 g14068(.a(new_n13958), .b(new_n13953), .O(new_n14262));
  inv1 g14069(.a(new_n14262), .O(new_n14263));
  nor2 g14070(.a(new_n14263), .b(new_n14261), .O(new_n14264));
  inv1 g14071(.a(new_n14261), .O(new_n14265));
  nor2 g14072(.a(new_n14262), .b(new_n14265), .O(new_n14266));
  nor2 g14073(.a(new_n14266), .b(new_n14264), .O(new_n14267));
  nor2 g14074(.a(new_n14065), .b(new_n14017), .O(new_n14268));
  inv1 g14075(.a(new_n14268), .O(new_n14269));
  nor2 g14076(.a(new_n14269), .b(new_n14267), .O(new_n14270));
  inv1 g14077(.a(new_n14267), .O(new_n14271));
  nor2 g14078(.a(new_n14268), .b(new_n14271), .O(new_n14272));
  nor2 g14079(.a(new_n14272), .b(new_n14270), .O(new_n14273));
  inv1 g14080(.a(new_n14273), .O(new_n14274));
  nor2 g14081(.a(new_n13982), .b(new_n13975), .O(new_n14275));
  nor2 g14082(.a(new_n14275), .b(new_n14274), .O(new_n14276));
  inv1 g14083(.a(new_n14275), .O(new_n14277));
  nor2 g14084(.a(new_n14277), .b(new_n14273), .O(new_n14278));
  nor2 g14085(.a(new_n14278), .b(new_n14276), .O(new_n14279));
  nor2 g14086(.a(new_n14279), .b(new_n14248), .O(new_n14280));
  inv1 g14087(.a(new_n14279), .O(new_n14281));
  nor2 g14088(.a(new_n14281), .b(new_n14247), .O(new_n14282));
  nor2 g14089(.a(new_n14282), .b(new_n14280), .O(new_n14283));
  nor2 g14090(.a(new_n14171), .b(new_n13985), .O(new_n14284));
  inv1 g14091(.a(new_n14284), .O(new_n14285));
  nor2 g14092(.a(new_n14285), .b(new_n14283), .O(new_n14286));
  inv1 g14093(.a(new_n14283), .O(new_n14287));
  nor2 g14094(.a(new_n14284), .b(new_n14287), .O(new_n14288));
  nor2 g14095(.a(new_n14288), .b(new_n14286), .O(new_n14289));
  nor2 g14096(.a(new_n14222), .b(new_n14216), .O(new_n14290));
  nor2 g14097(.a(new_n14162), .b(new_n14158), .O(new_n14291));
  nor2 g14098(.a(new_n14191), .b(new_n14185), .O(new_n14292));
  inv1 g14099(.a(new_n14292), .O(new_n14293));
  nor2 g14100(.a(new_n14062), .b(new_n14055), .O(new_n14294));
  inv1 g14101(.a(new_n14294), .O(new_n14295));
  nor2 g14102(.a(new_n14295), .b(new_n14293), .O(new_n14296));
  nor2 g14103(.a(new_n14294), .b(new_n14292), .O(new_n14297));
  nor2 g14104(.a(new_n14297), .b(new_n14296), .O(new_n14298));
  nor2 g14105(.a(new_n14155), .b(new_n14148), .O(new_n14299));
  inv1 g14106(.a(new_n14299), .O(new_n14300));
  nor2 g14107(.a(new_n14300), .b(new_n14298), .O(new_n14301));
  inv1 g14108(.a(new_n14298), .O(new_n14302));
  nor2 g14109(.a(new_n14299), .b(new_n14302), .O(new_n14303));
  nor2 g14110(.a(new_n14303), .b(new_n14301), .O(new_n14304));
  inv1 g14111(.a(new_n14304), .O(new_n14305));
  nor2 g14112(.a(new_n14305), .b(new_n14291), .O(new_n14306));
  inv1 g14113(.a(new_n14291), .O(new_n14307));
  nor2 g14114(.a(new_n14304), .b(new_n14307), .O(new_n14308));
  nor2 g14115(.a(new_n14308), .b(new_n14306), .O(new_n14309));
  inv1 g14116(.a(new_n14309), .O(new_n14310));
  nor2 g14117(.a(new_n14110), .b(new_n14104), .O(new_n14311));
  nor2 g14118(.a(new_n14030), .b(new_n14025), .O(new_n14312));
  nor2 g14119(.a(new_n14042), .b(new_n14035), .O(new_n14313));
  nor2 g14120(.a(new_n14313), .b(new_n14312), .O(new_n14314));
  inv1 g14121(.a(new_n14312), .O(new_n14315));
  inv1 g14122(.a(new_n14313), .O(new_n14316));
  nor2 g14123(.a(new_n14316), .b(new_n14315), .O(new_n14317));
  nor2 g14124(.a(new_n14317), .b(new_n14314), .O(new_n14318));
  nor2 g14125(.a(new_n14146), .b(new_n14139), .O(new_n14319));
  nor2 g14126(.a(new_n14319), .b(new_n14318), .O(new_n14320));
  inv1 g14127(.a(new_n14318), .O(new_n14321));
  inv1 g14128(.a(new_n14319), .O(new_n14322));
  nor2 g14129(.a(new_n14322), .b(new_n14321), .O(new_n14323));
  nor2 g14130(.a(new_n14323), .b(new_n14320), .O(new_n14324));
  nor2 g14131(.a(new_n14100), .b(new_n14097), .O(new_n14325));
  inv1 g14132(.a(new_n14325), .O(new_n14326));
  nor2 g14133(.a(new_n14088), .b(new_n14080), .O(new_n14327));
  nor2 g14134(.a(new_n14135), .b(new_n14129), .O(new_n14328));
  nor2 g14135(.a(new_n14328), .b(new_n14327), .O(new_n14329));
  inv1 g14136(.a(new_n14327), .O(new_n14330));
  inv1 g14137(.a(new_n14328), .O(new_n14331));
  nor2 g14138(.a(new_n14331), .b(new_n14330), .O(new_n14332));
  nor2 g14139(.a(new_n14332), .b(new_n14329), .O(new_n14333));
  nor2 g14140(.a(new_n14333), .b(new_n14326), .O(new_n14334));
  inv1 g14141(.a(new_n14333), .O(new_n14335));
  nor2 g14142(.a(new_n14335), .b(new_n14325), .O(new_n14336));
  nor2 g14143(.a(new_n14336), .b(new_n14334), .O(new_n14337));
  nor2 g14144(.a(new_n14337), .b(new_n14324), .O(new_n14338));
  inv1 g14145(.a(new_n14324), .O(new_n14339));
  inv1 g14146(.a(new_n14337), .O(new_n14340));
  nor2 g14147(.a(new_n14340), .b(new_n14339), .O(new_n14341));
  nor2 g14148(.a(new_n14341), .b(new_n14338), .O(new_n14342));
  inv1 g14149(.a(new_n14342), .O(new_n14343));
  nor2 g14150(.a(new_n14343), .b(new_n14311), .O(new_n14344));
  inv1 g14151(.a(new_n14311), .O(new_n14345));
  nor2 g14152(.a(new_n14342), .b(new_n14345), .O(new_n14346));
  nor2 g14153(.a(new_n14346), .b(new_n14344), .O(new_n14347));
  inv1 g14154(.a(new_n14347), .O(new_n14348));
  nor2 g14155(.a(new_n14348), .b(new_n14310), .O(new_n14349));
  nor2 g14156(.a(new_n14347), .b(new_n14309), .O(new_n14350));
  nor2 g14157(.a(new_n14350), .b(new_n14349), .O(new_n14351));
  inv1 g14158(.a(new_n14351), .O(new_n14352));
  nor2 g14159(.a(new_n14352), .b(new_n14290), .O(new_n14353));
  inv1 g14160(.a(new_n14290), .O(new_n14354));
  nor2 g14161(.a(new_n14351), .b(new_n14354), .O(new_n14355));
  nor2 g14162(.a(new_n14355), .b(new_n14353), .O(new_n14356));
  inv1 g14163(.a(new_n14356), .O(new_n14357));
  nor2 g14164(.a(new_n14211), .b(new_n14206), .O(new_n14358));
  nor2 g14165(.a(new_n14202), .b(new_n14199), .O(new_n14359));
  nor2 g14166(.a(new_n14053), .b(new_n14048), .O(new_n14360));
  nor2 g14167(.a(new_n14011), .b(new_n14003), .O(new_n14361));
  nor2 g14168(.a(new_n14361), .b(new_n14360), .O(new_n14362));
  inv1 g14169(.a(new_n14360), .O(new_n14363));
  inv1 g14170(.a(new_n14361), .O(new_n14364));
  nor2 g14171(.a(new_n14364), .b(new_n14363), .O(new_n14365));
  nor2 g14172(.a(new_n14365), .b(new_n14362), .O(new_n14366));
  inv1 g14173(.a(new_n14366), .O(new_n14367));
  nor2 g14174(.a(new_n11596), .b(new_n322), .O(new_n14368));
  nor2 g14175(.a(new_n10895), .b(new_n438), .O(new_n14369));
  nor2 g14176(.a(new_n14369), .b(new_n14368), .O(new_n14370));
  nor2 g14177(.a(new_n11596), .b(new_n438), .O(new_n14371));
  inv1 g14178(.a(new_n14371), .O(new_n14372));
  nor2 g14179(.a(new_n14372), .b(new_n13537), .O(new_n14373));
  nor2 g14180(.a(new_n14373), .b(new_n14370), .O(new_n14374));
  nor2 g14181(.a(new_n14374), .b(new_n14038), .O(new_n14375));
  inv1 g14182(.a(new_n14374), .O(new_n14376));
  nor2 g14183(.a(new_n14376), .b(new_n14037), .O(new_n14377));
  nor2 g14184(.a(new_n14377), .b(new_n14375), .O(new_n14378));
  nor2 g14185(.a(new_n14378), .b(new_n14367), .O(new_n14379));
  inv1 g14186(.a(new_n14378), .O(new_n14380));
  nor2 g14187(.a(new_n14380), .b(new_n14366), .O(new_n14381));
  nor2 g14188(.a(new_n14381), .b(new_n14379), .O(new_n14382));
  inv1 g14189(.a(new_n14382), .O(new_n14383));
  nor2 g14190(.a(new_n14383), .b(new_n14359), .O(new_n14384));
  inv1 g14191(.a(new_n14359), .O(new_n14385));
  nor2 g14192(.a(new_n14382), .b(new_n14385), .O(new_n14386));
  nor2 g14193(.a(new_n14386), .b(new_n14384), .O(new_n14387));
  inv1 g14194(.a(new_n14387), .O(new_n14388));
  nor2 g14195(.a(new_n7294), .b(new_n1425), .O(new_n14389));
  inv1 g14196(.a(new_n14389), .O(new_n14390));
  nor2 g14197(.a(new_n8026), .b(new_n1199), .O(new_n14391));
  nor2 g14198(.a(new_n14391), .b(new_n14118), .O(new_n14392));
  inv1 g14199(.a(new_n14115), .O(new_n14393));
  nor2 g14200(.a(new_n8026), .b(new_n1297), .O(new_n14394));
  inv1 g14201(.a(new_n14394), .O(new_n14395));
  nor2 g14202(.a(new_n14395), .b(new_n14393), .O(new_n14396));
  nor2 g14203(.a(new_n14396), .b(new_n14392), .O(new_n14397));
  nor2 g14204(.a(new_n14397), .b(new_n14390), .O(new_n14398));
  inv1 g14205(.a(new_n14397), .O(new_n14399));
  nor2 g14206(.a(new_n14399), .b(new_n14389), .O(new_n14400));
  nor2 g14207(.a(new_n14400), .b(new_n14398), .O(new_n14401));
  nor2 g14208(.a(new_n6958), .b(new_n1493), .O(new_n14402));
  inv1 g14209(.a(new_n14402), .O(new_n14403));
  nor2 g14210(.a(new_n11186), .b(new_n363), .O(new_n14404));
  nor2 g14211(.a(new_n14404), .b(\a[36] ), .O(new_n14405));
  nor2 g14212(.a(new_n11186), .b(new_n3870), .O(new_n14406));
  inv1 g14213(.a(new_n14406), .O(new_n14407));
  nor2 g14214(.a(new_n14407), .b(new_n363), .O(new_n14408));
  nor2 g14215(.a(new_n14408), .b(new_n14405), .O(new_n14409));
  nor2 g14216(.a(new_n14409), .b(new_n14403), .O(new_n14410));
  nor2 g14217(.a(new_n14405), .b(new_n14403), .O(new_n14411));
  nor2 g14218(.a(new_n14411), .b(new_n14408), .O(new_n14412));
  inv1 g14219(.a(new_n14412), .O(new_n14413));
  nor2 g14220(.a(new_n14413), .b(new_n14405), .O(new_n14414));
  nor2 g14221(.a(new_n14414), .b(new_n14410), .O(new_n14415));
  nor2 g14222(.a(new_n14415), .b(new_n14401), .O(new_n14416));
  inv1 g14223(.a(new_n14401), .O(new_n14417));
  inv1 g14224(.a(new_n14415), .O(new_n14418));
  nor2 g14225(.a(new_n14418), .b(new_n14417), .O(new_n14419));
  nor2 g14226(.a(new_n14419), .b(new_n14416), .O(new_n14420));
  inv1 g14227(.a(new_n14420), .O(new_n14421));
  nor2 g14228(.a(new_n4366), .b(new_n3231), .O(new_n14422));
  inv1 g14229(.a(new_n14422), .O(new_n14423));
  nor2 g14230(.a(new_n3870), .b(new_n3722), .O(new_n14424));
  nor2 g14231(.a(new_n14424), .b(new_n14005), .O(new_n14425));
  inv1 g14232(.a(new_n14424), .O(new_n14426));
  nor2 g14233(.a(new_n14426), .b(new_n14006), .O(new_n14427));
  nor2 g14234(.a(new_n14427), .b(new_n14425), .O(new_n14428));
  nor2 g14235(.a(new_n14428), .b(new_n14423), .O(new_n14429));
  inv1 g14236(.a(new_n14428), .O(new_n14430));
  nor2 g14237(.a(new_n14430), .b(new_n14422), .O(new_n14431));
  nor2 g14238(.a(new_n14431), .b(new_n14429), .O(new_n14432));
  nor2 g14239(.a(new_n14432), .b(new_n14421), .O(new_n14433));
  inv1 g14240(.a(new_n14432), .O(new_n14434));
  nor2 g14241(.a(new_n14434), .b(new_n14420), .O(new_n14435));
  nor2 g14242(.a(new_n14435), .b(new_n14433), .O(new_n14436));
  inv1 g14243(.a(new_n14436), .O(new_n14437));
  nor2 g14244(.a(new_n14437), .b(new_n14388), .O(new_n14438));
  nor2 g14245(.a(new_n14436), .b(new_n14387), .O(new_n14439));
  nor2 g14246(.a(new_n14439), .b(new_n14438), .O(new_n14440));
  inv1 g14247(.a(new_n14440), .O(new_n14441));
  nor2 g14248(.a(new_n14441), .b(new_n14358), .O(new_n14442));
  inv1 g14249(.a(new_n14358), .O(new_n14443));
  nor2 g14250(.a(new_n14440), .b(new_n14443), .O(new_n14444));
  nor2 g14251(.a(new_n14444), .b(new_n14442), .O(new_n14445));
  inv1 g14252(.a(new_n14445), .O(new_n14446));
  nor2 g14253(.a(new_n13972), .b(new_n13966), .O(new_n14447));
  nor2 g14254(.a(new_n9873), .b(new_n613), .O(new_n14448));
  nor2 g14255(.a(new_n10320), .b(new_n569), .O(new_n14449));
  nor2 g14256(.a(new_n14449), .b(new_n14448), .O(new_n14450));
  nor2 g14257(.a(new_n10320), .b(new_n613), .O(new_n14451));
  inv1 g14258(.a(new_n14451), .O(new_n14452));
  nor2 g14259(.a(new_n14452), .b(new_n14024), .O(new_n14453));
  nor2 g14260(.a(new_n14453), .b(new_n14450), .O(new_n14454));
  inv1 g14261(.a(new_n14454), .O(new_n14455));
  nor2 g14262(.a(new_n14124), .b(new_n14117), .O(new_n14456));
  inv1 g14263(.a(new_n14456), .O(new_n14457));
  nor2 g14264(.a(new_n14457), .b(new_n14455), .O(new_n14458));
  nor2 g14265(.a(new_n14456), .b(new_n14454), .O(new_n14459));
  nor2 g14266(.a(new_n14459), .b(new_n14458), .O(new_n14460));
  inv1 g14267(.a(new_n14460), .O(new_n14461));
  nor2 g14268(.a(new_n9658), .b(new_n699), .O(new_n14462));
  nor2 g14269(.a(new_n8946), .b(new_n847), .O(new_n14463));
  nor2 g14270(.a(new_n14463), .b(new_n14130), .O(new_n14464));
  inv1 g14271(.a(new_n14128), .O(new_n14465));
  nor2 g14272(.a(new_n14465), .b(new_n11980), .O(new_n14466));
  nor2 g14273(.a(new_n14466), .b(new_n14464), .O(new_n14467));
  inv1 g14274(.a(new_n14467), .O(new_n14468));
  nor2 g14275(.a(new_n14468), .b(new_n14462), .O(new_n14469));
  inv1 g14276(.a(new_n14462), .O(new_n14470));
  nor2 g14277(.a(new_n14467), .b(new_n14470), .O(new_n14471));
  nor2 g14278(.a(new_n14471), .b(new_n14469), .O(new_n14472));
  nor2 g14279(.a(new_n6570), .b(new_n1736), .O(new_n14473));
  inv1 g14280(.a(new_n14473), .O(new_n14474));
  nor2 g14281(.a(new_n6274), .b(new_n1903), .O(new_n14475));
  nor2 g14282(.a(new_n5971), .b(new_n2121), .O(new_n14476));
  nor2 g14283(.a(new_n14476), .b(new_n14475), .O(new_n14477));
  nor2 g14284(.a(new_n6274), .b(new_n2121), .O(new_n14478));
  inv1 g14285(.a(new_n14478), .O(new_n14479));
  nor2 g14286(.a(new_n14479), .b(new_n13746), .O(new_n14480));
  nor2 g14287(.a(new_n14480), .b(new_n14477), .O(new_n14481));
  nor2 g14288(.a(new_n14481), .b(new_n14474), .O(new_n14482));
  inv1 g14289(.a(new_n14481), .O(new_n14483));
  nor2 g14290(.a(new_n14483), .b(new_n14473), .O(new_n14484));
  nor2 g14291(.a(new_n14484), .b(new_n14482), .O(new_n14485));
  nor2 g14292(.a(new_n14485), .b(new_n14472), .O(new_n14486));
  inv1 g14293(.a(new_n14472), .O(new_n14487));
  inv1 g14294(.a(new_n14485), .O(new_n14488));
  nor2 g14295(.a(new_n14488), .b(new_n14487), .O(new_n14489));
  nor2 g14296(.a(new_n14489), .b(new_n14486), .O(new_n14490));
  inv1 g14297(.a(new_n14490), .O(new_n14491));
  nor2 g14298(.a(new_n14491), .b(new_n14461), .O(new_n14492));
  nor2 g14299(.a(new_n14490), .b(new_n14460), .O(new_n14493));
  nor2 g14300(.a(new_n14493), .b(new_n14492), .O(new_n14494));
  inv1 g14301(.a(new_n14494), .O(new_n14495));
  nor2 g14302(.a(new_n6893), .b(new_n1647), .O(new_n14496));
  inv1 g14303(.a(new_n14496), .O(new_n14497));
  nor2 g14304(.a(new_n8170), .b(new_n1086), .O(new_n14498));
  nor2 g14305(.a(new_n14498), .b(new_n11664), .O(new_n14499));
  inv1 g14306(.a(new_n14046), .O(new_n14500));
  nor2 g14307(.a(new_n14500), .b(new_n11287), .O(new_n14501));
  nor2 g14308(.a(new_n14501), .b(new_n14499), .O(new_n14502));
  nor2 g14309(.a(new_n14502), .b(new_n14497), .O(new_n14503));
  inv1 g14310(.a(new_n14502), .O(new_n14504));
  nor2 g14311(.a(new_n14504), .b(new_n14496), .O(new_n14505));
  nor2 g14312(.a(new_n14505), .b(new_n14503), .O(new_n14506));
  inv1 g14313(.a(new_n14506), .O(new_n14507));
  nor2 g14314(.a(new_n5393), .b(new_n2433), .O(new_n14508));
  nor2 g14315(.a(new_n5178), .b(new_n2506), .O(new_n14509));
  nor2 g14316(.a(new_n14509), .b(new_n14508), .O(new_n14510));
  nor2 g14317(.a(new_n5393), .b(new_n2506), .O(new_n14511));
  inv1 g14318(.a(new_n14511), .O(new_n14512));
  nor2 g14319(.a(new_n14512), .b(new_n14091), .O(new_n14513));
  nor2 g14320(.a(new_n14513), .b(new_n14510), .O(new_n14514));
  inv1 g14321(.a(new_n14514), .O(new_n14515));
  nor2 g14322(.a(new_n14515), .b(new_n14140), .O(new_n14516));
  nor2 g14323(.a(new_n14514), .b(new_n14141), .O(new_n14517));
  nor2 g14324(.a(new_n14517), .b(new_n14516), .O(new_n14518));
  nor2 g14325(.a(new_n4954), .b(new_n2660), .O(new_n14519));
  inv1 g14326(.a(new_n14519), .O(new_n14520));
  nor2 g14327(.a(new_n4425), .b(new_n3057), .O(new_n14521));
  nor2 g14328(.a(new_n14521), .b(new_n14082), .O(new_n14522));
  inv1 g14329(.a(new_n14079), .O(new_n14523));
  nor2 g14330(.a(new_n4682), .b(new_n3057), .O(new_n14524));
  inv1 g14331(.a(new_n14524), .O(new_n14525));
  nor2 g14332(.a(new_n14525), .b(new_n14523), .O(new_n14526));
  nor2 g14333(.a(new_n14526), .b(new_n14522), .O(new_n14527));
  nor2 g14334(.a(new_n14527), .b(new_n14520), .O(new_n14528));
  inv1 g14335(.a(new_n14527), .O(new_n14529));
  nor2 g14336(.a(new_n14529), .b(new_n14519), .O(new_n14530));
  nor2 g14337(.a(new_n14530), .b(new_n14528), .O(new_n14531));
  nor2 g14338(.a(new_n14531), .b(new_n14518), .O(new_n14532));
  inv1 g14339(.a(new_n14518), .O(new_n14533));
  inv1 g14340(.a(new_n14531), .O(new_n14534));
  nor2 g14341(.a(new_n14534), .b(new_n14533), .O(new_n14535));
  nor2 g14342(.a(new_n14535), .b(new_n14532), .O(new_n14536));
  nor2 g14343(.a(new_n14536), .b(new_n14507), .O(new_n14537));
  inv1 g14344(.a(new_n14536), .O(new_n14538));
  nor2 g14345(.a(new_n14538), .b(new_n14506), .O(new_n14539));
  nor2 g14346(.a(new_n14539), .b(new_n14537), .O(new_n14540));
  inv1 g14347(.a(new_n14540), .O(new_n14541));
  nor2 g14348(.a(new_n14541), .b(new_n14495), .O(new_n14542));
  nor2 g14349(.a(new_n14540), .b(new_n14494), .O(new_n14543));
  nor2 g14350(.a(new_n14543), .b(new_n14542), .O(new_n14544));
  inv1 g14351(.a(new_n14544), .O(new_n14545));
  nor2 g14352(.a(new_n14545), .b(new_n14447), .O(new_n14546));
  inv1 g14353(.a(new_n14447), .O(new_n14547));
  nor2 g14354(.a(new_n14544), .b(new_n14547), .O(new_n14548));
  nor2 g14355(.a(new_n14548), .b(new_n14546), .O(new_n14549));
  inv1 g14356(.a(new_n14549), .O(new_n14550));
  nor2 g14357(.a(new_n14550), .b(new_n14446), .O(new_n14551));
  nor2 g14358(.a(new_n14549), .b(new_n14445), .O(new_n14552));
  nor2 g14359(.a(new_n14552), .b(new_n14551), .O(new_n14553));
  inv1 g14360(.a(new_n14553), .O(new_n14554));
  nor2 g14361(.a(new_n14554), .b(new_n14357), .O(new_n14555));
  nor2 g14362(.a(new_n14553), .b(new_n14356), .O(new_n14556));
  nor2 g14363(.a(new_n14556), .b(new_n14555), .O(new_n14557));
  nor2 g14364(.a(new_n14557), .b(new_n14289), .O(new_n14558));
  inv1 g14365(.a(new_n14289), .O(new_n14559));
  inv1 g14366(.a(new_n14557), .O(new_n14560));
  nor2 g14367(.a(new_n14560), .b(new_n14559), .O(new_n14561));
  nor2 g14368(.a(new_n14561), .b(new_n14558), .O(new_n14562));
  nor2 g14369(.a(new_n14562), .b(new_n14246), .O(new_n14563));
  inv1 g14370(.a(new_n14562), .O(new_n14564));
  nor2 g14371(.a(new_n14564), .b(new_n14245), .O(new_n14565));
  nor2 g14372(.a(new_n14565), .b(new_n14563), .O(new_n14566));
  inv1 g14373(.a(new_n14566), .O(new_n14567));
  nor2 g14374(.a(new_n14240), .b(new_n14234), .O(new_n14568));
  nor2 g14375(.a(new_n14568), .b(new_n14567), .O(new_n14569));
  inv1 g14376(.a(new_n14568), .O(new_n14570));
  nor2 g14377(.a(new_n14570), .b(new_n14566), .O(new_n14571));
  nor2 g14378(.a(new_n14571), .b(new_n14569), .O(new_n14572));
  inv1 g14379(.a(new_n14572), .O(\asquared[72] ));
  nor2 g14380(.a(new_n14551), .b(new_n14442), .O(new_n14574));
  inv1 g14381(.a(new_n14574), .O(new_n14575));
  nor2 g14382(.a(new_n14344), .b(new_n14341), .O(new_n14576));
  nor2 g14383(.a(new_n14336), .b(new_n14332), .O(new_n14577));
  inv1 g14384(.a(new_n14577), .O(new_n14578));
  nor2 g14385(.a(new_n4954), .b(new_n2826), .O(new_n14579));
  nor2 g14386(.a(new_n5178), .b(new_n2660), .O(new_n14580));
  nor2 g14387(.a(new_n14580), .b(new_n14579), .O(new_n14581));
  nor2 g14388(.a(new_n5178), .b(new_n2826), .O(new_n14582));
  inv1 g14389(.a(new_n14582), .O(new_n14583));
  nor2 g14390(.a(new_n14583), .b(new_n14520), .O(new_n14584));
  nor2 g14391(.a(new_n14584), .b(new_n14581), .O(new_n14585));
  nor2 g14392(.a(new_n14585), .b(new_n14512), .O(new_n14586));
  inv1 g14393(.a(new_n14585), .O(new_n14587));
  nor2 g14394(.a(new_n14587), .b(new_n14511), .O(new_n14588));
  nor2 g14395(.a(new_n14588), .b(new_n14586), .O(new_n14589));
  nor2 g14396(.a(new_n14379), .b(new_n14365), .O(new_n14590));
  nor2 g14397(.a(new_n14590), .b(new_n14589), .O(new_n14591));
  inv1 g14398(.a(new_n14589), .O(new_n14592));
  inv1 g14399(.a(new_n14590), .O(new_n14593));
  nor2 g14400(.a(new_n14593), .b(new_n14592), .O(new_n14594));
  nor2 g14401(.a(new_n14594), .b(new_n14591), .O(new_n14595));
  nor2 g14402(.a(new_n14595), .b(new_n14578), .O(new_n14596));
  inv1 g14403(.a(new_n14595), .O(new_n14597));
  nor2 g14404(.a(new_n14597), .b(new_n14577), .O(new_n14598));
  nor2 g14405(.a(new_n14598), .b(new_n14596), .O(new_n14599));
  inv1 g14406(.a(new_n14599), .O(new_n14600));
  nor2 g14407(.a(new_n14600), .b(new_n14576), .O(new_n14601));
  inv1 g14408(.a(new_n14576), .O(new_n14602));
  nor2 g14409(.a(new_n14599), .b(new_n14602), .O(new_n14603));
  nor2 g14410(.a(new_n14603), .b(new_n14601), .O(new_n14604));
  nor2 g14411(.a(new_n14438), .b(new_n14384), .O(new_n14605));
  inv1 g14412(.a(new_n14605), .O(new_n14606));
  nor2 g14413(.a(new_n14606), .b(new_n14604), .O(new_n14607));
  inv1 g14414(.a(new_n14604), .O(new_n14608));
  nor2 g14415(.a(new_n14605), .b(new_n14608), .O(new_n14609));
  nor2 g14416(.a(new_n14609), .b(new_n14607), .O(new_n14610));
  inv1 g14417(.a(new_n14610), .O(new_n14611));
  nor2 g14418(.a(new_n14349), .b(new_n14306), .O(new_n14612));
  nor2 g14419(.a(new_n14612), .b(new_n14611), .O(new_n14613));
  inv1 g14420(.a(new_n14612), .O(new_n14614));
  nor2 g14421(.a(new_n14614), .b(new_n14610), .O(new_n14615));
  nor2 g14422(.a(new_n14615), .b(new_n14613), .O(new_n14616));
  nor2 g14423(.a(new_n14616), .b(new_n14575), .O(new_n14617));
  inv1 g14424(.a(new_n14616), .O(new_n14618));
  nor2 g14425(.a(new_n14618), .b(new_n14574), .O(new_n14619));
  nor2 g14426(.a(new_n14619), .b(new_n14617), .O(new_n14620));
  nor2 g14427(.a(new_n14555), .b(new_n14353), .O(new_n14621));
  inv1 g14428(.a(new_n14621), .O(new_n14622));
  nor2 g14429(.a(new_n14622), .b(new_n14620), .O(new_n14623));
  inv1 g14430(.a(new_n14620), .O(new_n14624));
  nor2 g14431(.a(new_n14621), .b(new_n14624), .O(new_n14625));
  nor2 g14432(.a(new_n14625), .b(new_n14623), .O(new_n14626));
  nor2 g14433(.a(new_n14282), .b(new_n14276), .O(new_n14627));
  inv1 g14434(.a(new_n14627), .O(new_n14628));
  nor2 g14435(.a(new_n14323), .b(new_n14317), .O(new_n14629));
  inv1 g14436(.a(new_n14629), .O(new_n14630));
  nor2 g14437(.a(new_n14539), .b(new_n14532), .O(new_n14631));
  inv1 g14438(.a(new_n14631), .O(new_n14632));
  nor2 g14439(.a(new_n14632), .b(new_n14630), .O(new_n14633));
  nor2 g14440(.a(new_n14631), .b(new_n14629), .O(new_n14634));
  nor2 g14441(.a(new_n14634), .b(new_n14633), .O(new_n14635));
  nor2 g14442(.a(new_n14433), .b(new_n14416), .O(new_n14636));
  inv1 g14443(.a(new_n14636), .O(new_n14637));
  nor2 g14444(.a(new_n14637), .b(new_n14635), .O(new_n14638));
  inv1 g14445(.a(new_n14635), .O(new_n14639));
  nor2 g14446(.a(new_n14636), .b(new_n14639), .O(new_n14640));
  nor2 g14447(.a(new_n14640), .b(new_n14638), .O(new_n14641));
  nor2 g14448(.a(new_n14546), .b(new_n14542), .O(new_n14642));
  inv1 g14449(.a(new_n14642), .O(new_n14643));
  nor2 g14450(.a(new_n14643), .b(new_n14641), .O(new_n14644));
  inv1 g14451(.a(new_n14641), .O(new_n14645));
  nor2 g14452(.a(new_n14642), .b(new_n14645), .O(new_n14646));
  nor2 g14453(.a(new_n14646), .b(new_n14644), .O(new_n14647));
  inv1 g14454(.a(new_n14647), .O(new_n14648));
  nor2 g14455(.a(new_n14492), .b(new_n14486), .O(new_n14649));
  nor2 g14456(.a(new_n14505), .b(new_n14499), .O(new_n14650));
  nor2 g14457(.a(new_n14516), .b(new_n14510), .O(new_n14651));
  nor2 g14458(.a(new_n14651), .b(new_n14650), .O(new_n14652));
  inv1 g14459(.a(new_n14650), .O(new_n14653));
  inv1 g14460(.a(new_n14651), .O(new_n14654));
  nor2 g14461(.a(new_n14654), .b(new_n14653), .O(new_n14655));
  nor2 g14462(.a(new_n14655), .b(new_n14652), .O(new_n14656));
  nor2 g14463(.a(new_n14530), .b(new_n14522), .O(new_n14657));
  nor2 g14464(.a(new_n14657), .b(new_n14656), .O(new_n14658));
  inv1 g14465(.a(new_n14656), .O(new_n14659));
  inv1 g14466(.a(new_n14657), .O(new_n14660));
  nor2 g14467(.a(new_n14660), .b(new_n14659), .O(new_n14661));
  nor2 g14468(.a(new_n14661), .b(new_n14658), .O(new_n14662));
  inv1 g14469(.a(new_n14662), .O(new_n14663));
  nor2 g14470(.a(new_n14431), .b(new_n14425), .O(new_n14664));
  nor2 g14471(.a(new_n14664), .b(new_n14413), .O(new_n14665));
  inv1 g14472(.a(new_n14664), .O(new_n14666));
  nor2 g14473(.a(new_n14666), .b(new_n14412), .O(new_n14667));
  nor2 g14474(.a(new_n14667), .b(new_n14665), .O(new_n14668));
  nor2 g14475(.a(new_n14400), .b(new_n14392), .O(new_n14669));
  nor2 g14476(.a(new_n14669), .b(new_n14668), .O(new_n14670));
  inv1 g14477(.a(new_n14668), .O(new_n14671));
  inv1 g14478(.a(new_n14669), .O(new_n14672));
  nor2 g14479(.a(new_n14672), .b(new_n14671), .O(new_n14673));
  nor2 g14480(.a(new_n14673), .b(new_n14670), .O(new_n14674));
  inv1 g14481(.a(new_n14674), .O(new_n14675));
  nor2 g14482(.a(new_n14675), .b(new_n14663), .O(new_n14676));
  nor2 g14483(.a(new_n14674), .b(new_n14662), .O(new_n14677));
  nor2 g14484(.a(new_n14677), .b(new_n14676), .O(new_n14678));
  inv1 g14485(.a(new_n14678), .O(new_n14679));
  nor2 g14486(.a(new_n14679), .b(new_n14649), .O(new_n14680));
  inv1 g14487(.a(new_n14649), .O(new_n14681));
  nor2 g14488(.a(new_n14678), .b(new_n14681), .O(new_n14682));
  nor2 g14489(.a(new_n14682), .b(new_n14680), .O(new_n14683));
  inv1 g14490(.a(new_n14683), .O(new_n14684));
  nor2 g14491(.a(new_n14684), .b(new_n14648), .O(new_n14685));
  nor2 g14492(.a(new_n14683), .b(new_n14647), .O(new_n14686));
  nor2 g14493(.a(new_n14686), .b(new_n14685), .O(new_n14687));
  nor2 g14494(.a(new_n14687), .b(new_n14628), .O(new_n14688));
  inv1 g14495(.a(new_n14687), .O(new_n14689));
  nor2 g14496(.a(new_n14689), .b(new_n14627), .O(new_n14690));
  nor2 g14497(.a(new_n14690), .b(new_n14688), .O(new_n14691));
  inv1 g14498(.a(new_n14691), .O(new_n14692));
  nor2 g14499(.a(new_n14303), .b(new_n14297), .O(new_n14693));
  nor2 g14500(.a(new_n11596), .b(new_n363), .O(new_n14694));
  nor2 g14501(.a(new_n11186), .b(new_n438), .O(new_n14695));
  nor2 g14502(.a(new_n10895), .b(new_n502), .O(new_n14696));
  nor2 g14503(.a(new_n14696), .b(new_n14695), .O(new_n14697));
  inv1 g14504(.a(new_n14369), .O(new_n14698));
  nor2 g14505(.a(new_n11186), .b(new_n502), .O(new_n14699));
  inv1 g14506(.a(new_n14699), .O(new_n14700));
  nor2 g14507(.a(new_n14700), .b(new_n14698), .O(new_n14701));
  nor2 g14508(.a(new_n14701), .b(new_n14697), .O(new_n14702));
  inv1 g14509(.a(new_n14702), .O(new_n14703));
  nor2 g14510(.a(new_n14703), .b(new_n14694), .O(new_n14704));
  inv1 g14511(.a(new_n14694), .O(new_n14705));
  nor2 g14512(.a(new_n14702), .b(new_n14705), .O(new_n14706));
  nor2 g14513(.a(new_n14706), .b(new_n14704), .O(new_n14707));
  nor2 g14514(.a(new_n14458), .b(new_n14453), .O(new_n14708));
  nor2 g14515(.a(new_n10468), .b(new_n569), .O(new_n14709));
  inv1 g14516(.a(new_n14709), .O(new_n14710));
  nor2 g14517(.a(new_n6893), .b(new_n1736), .O(new_n14711));
  nor2 g14518(.a(new_n6570), .b(new_n1903), .O(new_n14712));
  nor2 g14519(.a(new_n14712), .b(new_n14711), .O(new_n14713));
  nor2 g14520(.a(new_n6893), .b(new_n1903), .O(new_n14714));
  inv1 g14521(.a(new_n14714), .O(new_n14715));
  nor2 g14522(.a(new_n14715), .b(new_n14474), .O(new_n14716));
  nor2 g14523(.a(new_n14716), .b(new_n14713), .O(new_n14717));
  nor2 g14524(.a(new_n14717), .b(new_n14710), .O(new_n14718));
  inv1 g14525(.a(new_n14717), .O(new_n14719));
  nor2 g14526(.a(new_n14719), .b(new_n14709), .O(new_n14720));
  nor2 g14527(.a(new_n14720), .b(new_n14718), .O(new_n14721));
  nor2 g14528(.a(new_n14721), .b(new_n14708), .O(new_n14722));
  inv1 g14529(.a(new_n14708), .O(new_n14723));
  inv1 g14530(.a(new_n14721), .O(new_n14724));
  nor2 g14531(.a(new_n14724), .b(new_n14723), .O(new_n14725));
  nor2 g14532(.a(new_n14725), .b(new_n14722), .O(new_n14726));
  inv1 g14533(.a(new_n14726), .O(new_n14727));
  nor2 g14534(.a(new_n14727), .b(new_n14707), .O(new_n14728));
  inv1 g14535(.a(new_n14707), .O(new_n14729));
  nor2 g14536(.a(new_n14726), .b(new_n14729), .O(new_n14730));
  nor2 g14537(.a(new_n14730), .b(new_n14728), .O(new_n14731));
  inv1 g14538(.a(new_n14731), .O(new_n14732));
  nor2 g14539(.a(new_n4093), .b(new_n3722), .O(new_n14733));
  inv1 g14540(.a(new_n14733), .O(new_n14734));
  nor2 g14541(.a(new_n7537), .b(new_n1425), .O(new_n14735));
  nor2 g14542(.a(new_n7294), .b(new_n1493), .O(new_n14736));
  nor2 g14543(.a(new_n14736), .b(new_n14735), .O(new_n14737));
  nor2 g14544(.a(new_n7537), .b(new_n1493), .O(new_n14738));
  inv1 g14545(.a(new_n14738), .O(new_n14739));
  nor2 g14546(.a(new_n14739), .b(new_n14390), .O(new_n14740));
  nor2 g14547(.a(new_n14740), .b(new_n14737), .O(new_n14741));
  nor2 g14548(.a(new_n14741), .b(new_n14734), .O(new_n14742));
  inv1 g14549(.a(new_n14741), .O(new_n14743));
  nor2 g14550(.a(new_n14743), .b(new_n14733), .O(new_n14744));
  nor2 g14551(.a(new_n14744), .b(new_n14742), .O(new_n14745));
  nor2 g14552(.a(new_n6958), .b(new_n1647), .O(new_n14746));
  nor2 g14553(.a(new_n14746), .b(new_n11979), .O(new_n14747));
  inv1 g14554(.a(new_n14746), .O(new_n14748));
  nor2 g14555(.a(new_n14748), .b(new_n11980), .O(new_n14749));
  nor2 g14556(.a(new_n14749), .b(new_n14747), .O(new_n14750));
  inv1 g14557(.a(new_n14750), .O(new_n14751));
  nor2 g14558(.a(new_n14751), .b(new_n14525), .O(new_n14752));
  nor2 g14559(.a(new_n14750), .b(new_n14524), .O(new_n14753));
  nor2 g14560(.a(new_n14753), .b(new_n14752), .O(new_n14754));
  inv1 g14561(.a(new_n14754), .O(new_n14755));
  nor2 g14562(.a(new_n14755), .b(new_n14745), .O(new_n14756));
  inv1 g14563(.a(new_n14745), .O(new_n14757));
  nor2 g14564(.a(new_n14754), .b(new_n14757), .O(new_n14758));
  nor2 g14565(.a(new_n14758), .b(new_n14756), .O(new_n14759));
  inv1 g14566(.a(new_n14759), .O(new_n14760));
  nor2 g14567(.a(new_n8946), .b(new_n941), .O(new_n14761));
  inv1 g14568(.a(new_n14761), .O(new_n14762));
  nor2 g14569(.a(new_n14394), .b(new_n11286), .O(new_n14763));
  nor2 g14570(.a(new_n8476), .b(new_n1297), .O(new_n14764));
  inv1 g14571(.a(new_n14764), .O(new_n14765));
  nor2 g14572(.a(new_n14765), .b(new_n10280), .O(new_n14766));
  nor2 g14573(.a(new_n14766), .b(new_n14763), .O(new_n14767));
  nor2 g14574(.a(new_n14767), .b(new_n14762), .O(new_n14768));
  inv1 g14575(.a(new_n14767), .O(new_n14769));
  nor2 g14576(.a(new_n14769), .b(new_n14761), .O(new_n14770));
  nor2 g14577(.a(new_n14770), .b(new_n14768), .O(new_n14771));
  nor2 g14578(.a(new_n14771), .b(new_n14760), .O(new_n14772));
  inv1 g14579(.a(new_n14771), .O(new_n14773));
  nor2 g14580(.a(new_n14773), .b(new_n14759), .O(new_n14774));
  nor2 g14581(.a(new_n14774), .b(new_n14772), .O(new_n14775));
  inv1 g14582(.a(new_n14775), .O(new_n14776));
  nor2 g14583(.a(new_n14776), .b(new_n14732), .O(new_n14777));
  nor2 g14584(.a(new_n14775), .b(new_n14731), .O(new_n14778));
  nor2 g14585(.a(new_n14778), .b(new_n14777), .O(new_n14779));
  inv1 g14586(.a(new_n14779), .O(new_n14780));
  nor2 g14587(.a(new_n14780), .b(new_n14693), .O(new_n14781));
  inv1 g14588(.a(new_n14693), .O(new_n14782));
  nor2 g14589(.a(new_n14779), .b(new_n14782), .O(new_n14783));
  nor2 g14590(.a(new_n14783), .b(new_n14781), .O(new_n14784));
  inv1 g14591(.a(new_n14784), .O(new_n14785));
  nor2 g14592(.a(new_n14272), .b(new_n14266), .O(new_n14786));
  nor2 g14593(.a(new_n14484), .b(new_n14477), .O(new_n14787));
  nor2 g14594(.a(new_n14469), .b(new_n14464), .O(new_n14788));
  nor2 g14595(.a(new_n14788), .b(new_n14787), .O(new_n14789));
  inv1 g14596(.a(new_n14787), .O(new_n14790));
  inv1 g14597(.a(new_n14788), .O(new_n14791));
  nor2 g14598(.a(new_n14791), .b(new_n14790), .O(new_n14792));
  nor2 g14599(.a(new_n14792), .b(new_n14789), .O(new_n14793));
  nor2 g14600(.a(new_n14377), .b(new_n14370), .O(new_n14794));
  nor2 g14601(.a(new_n14794), .b(new_n14793), .O(new_n14795));
  inv1 g14602(.a(new_n14793), .O(new_n14796));
  inv1 g14603(.a(new_n14794), .O(new_n14797));
  nor2 g14604(.a(new_n14797), .b(new_n14796), .O(new_n14798));
  nor2 g14605(.a(new_n14798), .b(new_n14795), .O(new_n14799));
  nor2 g14606(.a(new_n14260), .b(new_n14254), .O(new_n14800));
  inv1 g14607(.a(new_n14800), .O(new_n14801));
  nor2 g14608(.a(new_n14801), .b(new_n14799), .O(new_n14802));
  inv1 g14609(.a(new_n14799), .O(new_n14803));
  nor2 g14610(.a(new_n14800), .b(new_n14803), .O(new_n14804));
  nor2 g14611(.a(new_n14804), .b(new_n14802), .O(new_n14805));
  nor2 g14612(.a(new_n8170), .b(new_n1199), .O(new_n14806));
  inv1 g14613(.a(new_n14806), .O(new_n14807));
  nor2 g14614(.a(new_n4366), .b(new_n3533), .O(new_n14808));
  nor2 g14615(.a(new_n4425), .b(new_n3231), .O(new_n14809));
  nor2 g14616(.a(new_n14809), .b(new_n14808), .O(new_n14810));
  nor2 g14617(.a(new_n4425), .b(new_n3533), .O(new_n14811));
  inv1 g14618(.a(new_n14811), .O(new_n14812));
  nor2 g14619(.a(new_n14812), .b(new_n14423), .O(new_n14813));
  nor2 g14620(.a(new_n14813), .b(new_n14810), .O(new_n14814));
  nor2 g14621(.a(new_n14814), .b(new_n14807), .O(new_n14815));
  inv1 g14622(.a(new_n14814), .O(new_n14816));
  nor2 g14623(.a(new_n14816), .b(new_n14806), .O(new_n14817));
  nor2 g14624(.a(new_n14817), .b(new_n14815), .O(new_n14818));
  inv1 g14625(.a(new_n14818), .O(new_n14819));
  nor2 g14626(.a(new_n9873), .b(new_n699), .O(new_n14820));
  nor2 g14627(.a(new_n9658), .b(new_n800), .O(new_n14821));
  nor2 g14628(.a(new_n14821), .b(new_n14820), .O(new_n14822));
  nor2 g14629(.a(new_n9873), .b(new_n800), .O(new_n14823));
  inv1 g14630(.a(new_n14823), .O(new_n14824));
  nor2 g14631(.a(new_n14824), .b(new_n14470), .O(new_n14825));
  nor2 g14632(.a(new_n14825), .b(new_n14822), .O(new_n14826));
  inv1 g14633(.a(new_n14826), .O(new_n14827));
  nor2 g14634(.a(new_n14827), .b(new_n14451), .O(new_n14828));
  nor2 g14635(.a(new_n14826), .b(new_n14452), .O(new_n14829));
  nor2 g14636(.a(new_n14829), .b(new_n14828), .O(new_n14830));
  nor2 g14637(.a(new_n5971), .b(new_n2184), .O(new_n14831));
  nor2 g14638(.a(new_n5796), .b(new_n2433), .O(new_n14832));
  nor2 g14639(.a(new_n14832), .b(new_n14831), .O(new_n14833));
  nor2 g14640(.a(new_n5971), .b(new_n2433), .O(new_n14834));
  inv1 g14641(.a(new_n14834), .O(new_n14835));
  nor2 g14642(.a(new_n14835), .b(new_n14141), .O(new_n14836));
  nor2 g14643(.a(new_n14836), .b(new_n14833), .O(new_n14837));
  nor2 g14644(.a(new_n14837), .b(new_n14479), .O(new_n14838));
  inv1 g14645(.a(new_n14837), .O(new_n14839));
  nor2 g14646(.a(new_n14839), .b(new_n14478), .O(new_n14840));
  nor2 g14647(.a(new_n14840), .b(new_n14838), .O(new_n14841));
  nor2 g14648(.a(new_n14841), .b(new_n14830), .O(new_n14842));
  inv1 g14649(.a(new_n14830), .O(new_n14843));
  inv1 g14650(.a(new_n14841), .O(new_n14844));
  nor2 g14651(.a(new_n14844), .b(new_n14843), .O(new_n14845));
  nor2 g14652(.a(new_n14845), .b(new_n14842), .O(new_n14846));
  nor2 g14653(.a(new_n14846), .b(new_n14819), .O(new_n14847));
  inv1 g14654(.a(new_n14846), .O(new_n14848));
  nor2 g14655(.a(new_n14848), .b(new_n14818), .O(new_n14849));
  nor2 g14656(.a(new_n14849), .b(new_n14847), .O(new_n14850));
  nor2 g14657(.a(new_n14850), .b(new_n14805), .O(new_n14851));
  inv1 g14658(.a(new_n14805), .O(new_n14852));
  inv1 g14659(.a(new_n14850), .O(new_n14853));
  nor2 g14660(.a(new_n14853), .b(new_n14852), .O(new_n14854));
  nor2 g14661(.a(new_n14854), .b(new_n14851), .O(new_n14855));
  inv1 g14662(.a(new_n14855), .O(new_n14856));
  nor2 g14663(.a(new_n14856), .b(new_n14786), .O(new_n14857));
  inv1 g14664(.a(new_n14786), .O(new_n14858));
  nor2 g14665(.a(new_n14855), .b(new_n14858), .O(new_n14859));
  nor2 g14666(.a(new_n14859), .b(new_n14857), .O(new_n14860));
  inv1 g14667(.a(new_n14860), .O(new_n14861));
  nor2 g14668(.a(new_n14861), .b(new_n14785), .O(new_n14862));
  nor2 g14669(.a(new_n14860), .b(new_n14784), .O(new_n14863));
  nor2 g14670(.a(new_n14863), .b(new_n14862), .O(new_n14864));
  inv1 g14671(.a(new_n14864), .O(new_n14865));
  nor2 g14672(.a(new_n14865), .b(new_n14692), .O(new_n14866));
  nor2 g14673(.a(new_n14864), .b(new_n14691), .O(new_n14867));
  nor2 g14674(.a(new_n14867), .b(new_n14866), .O(new_n14868));
  nor2 g14675(.a(new_n14868), .b(new_n14626), .O(new_n14869));
  inv1 g14676(.a(new_n14626), .O(new_n14870));
  inv1 g14677(.a(new_n14868), .O(new_n14871));
  nor2 g14678(.a(new_n14871), .b(new_n14870), .O(new_n14872));
  nor2 g14679(.a(new_n14872), .b(new_n14869), .O(new_n14873));
  nor2 g14680(.a(new_n14561), .b(new_n14288), .O(new_n14874));
  inv1 g14681(.a(new_n14874), .O(new_n14875));
  nor2 g14682(.a(new_n14875), .b(new_n14873), .O(new_n14876));
  inv1 g14683(.a(new_n14873), .O(new_n14877));
  nor2 g14684(.a(new_n14874), .b(new_n14877), .O(new_n14878));
  nor2 g14685(.a(new_n14878), .b(new_n14876), .O(new_n14879));
  nor2 g14686(.a(new_n14569), .b(new_n14563), .O(new_n14880));
  inv1 g14687(.a(new_n14880), .O(new_n14881));
  nor2 g14688(.a(new_n14881), .b(new_n14879), .O(new_n14882));
  inv1 g14689(.a(new_n14879), .O(new_n14883));
  nor2 g14690(.a(new_n14880), .b(new_n14883), .O(new_n14884));
  nor2 g14691(.a(new_n14884), .b(new_n14882), .O(new_n14885));
  inv1 g14692(.a(new_n14885), .O(\asquared[73] ));
  nor2 g14693(.a(new_n14872), .b(new_n14625), .O(new_n14887));
  inv1 g14694(.a(new_n14887), .O(new_n14888));
  nor2 g14695(.a(new_n14866), .b(new_n14690), .O(new_n14889));
  inv1 g14696(.a(new_n14889), .O(new_n14890));
  nor2 g14697(.a(new_n14862), .b(new_n14857), .O(new_n14891));
  nor2 g14698(.a(new_n14685), .b(new_n14646), .O(new_n14892));
  nor2 g14699(.a(new_n14854), .b(new_n14804), .O(new_n14893));
  nor2 g14700(.a(new_n14661), .b(new_n14655), .O(new_n14894));
  inv1 g14701(.a(new_n14894), .O(new_n14895));
  nor2 g14702(.a(new_n14798), .b(new_n14792), .O(new_n14896));
  nor2 g14703(.a(new_n4954), .b(new_n3057), .O(new_n14897));
  nor2 g14704(.a(new_n4682), .b(new_n3231), .O(new_n14898));
  nor2 g14705(.a(new_n14898), .b(new_n14897), .O(new_n14899));
  nor2 g14706(.a(new_n4954), .b(new_n3231), .O(new_n14900));
  inv1 g14707(.a(new_n14900), .O(new_n14901));
  nor2 g14708(.a(new_n14901), .b(new_n14525), .O(new_n14902));
  nor2 g14709(.a(new_n14902), .b(new_n14899), .O(new_n14903));
  nor2 g14710(.a(new_n14903), .b(new_n14583), .O(new_n14904));
  inv1 g14711(.a(new_n14903), .O(new_n14905));
  nor2 g14712(.a(new_n14905), .b(new_n14582), .O(new_n14906));
  nor2 g14713(.a(new_n14906), .b(new_n14904), .O(new_n14907));
  nor2 g14714(.a(new_n14907), .b(new_n14896), .O(new_n14908));
  inv1 g14715(.a(new_n14896), .O(new_n14909));
  inv1 g14716(.a(new_n14907), .O(new_n14910));
  nor2 g14717(.a(new_n14910), .b(new_n14909), .O(new_n14911));
  nor2 g14718(.a(new_n14911), .b(new_n14908), .O(new_n14912));
  nor2 g14719(.a(new_n14912), .b(new_n14895), .O(new_n14913));
  inv1 g14720(.a(new_n14912), .O(new_n14914));
  nor2 g14721(.a(new_n14914), .b(new_n14894), .O(new_n14915));
  nor2 g14722(.a(new_n14915), .b(new_n14913), .O(new_n14916));
  inv1 g14723(.a(new_n14916), .O(new_n14917));
  nor2 g14724(.a(new_n14680), .b(new_n14676), .O(new_n14918));
  nor2 g14725(.a(new_n14918), .b(new_n14917), .O(new_n14919));
  inv1 g14726(.a(new_n14918), .O(new_n14920));
  nor2 g14727(.a(new_n14920), .b(new_n14916), .O(new_n14921));
  nor2 g14728(.a(new_n14921), .b(new_n14919), .O(new_n14922));
  inv1 g14729(.a(new_n14922), .O(new_n14923));
  nor2 g14730(.a(new_n14923), .b(new_n14893), .O(new_n14924));
  inv1 g14731(.a(new_n14893), .O(new_n14925));
  nor2 g14732(.a(new_n14922), .b(new_n14925), .O(new_n14926));
  nor2 g14733(.a(new_n14926), .b(new_n14924), .O(new_n14927));
  inv1 g14734(.a(new_n14927), .O(new_n14928));
  nor2 g14735(.a(new_n14928), .b(new_n14892), .O(new_n14929));
  inv1 g14736(.a(new_n14892), .O(new_n14930));
  nor2 g14737(.a(new_n14927), .b(new_n14930), .O(new_n14931));
  nor2 g14738(.a(new_n14931), .b(new_n14929), .O(new_n14932));
  inv1 g14739(.a(new_n14932), .O(new_n14933));
  nor2 g14740(.a(new_n14933), .b(new_n14891), .O(new_n14934));
  inv1 g14741(.a(new_n14891), .O(new_n14935));
  nor2 g14742(.a(new_n14932), .b(new_n14935), .O(new_n14936));
  nor2 g14743(.a(new_n14936), .b(new_n14934), .O(new_n14937));
  nor2 g14744(.a(new_n14937), .b(new_n14890), .O(new_n14938));
  inv1 g14745(.a(new_n14937), .O(new_n14939));
  nor2 g14746(.a(new_n14939), .b(new_n14889), .O(new_n14940));
  nor2 g14747(.a(new_n14940), .b(new_n14938), .O(new_n14941));
  nor2 g14748(.a(new_n14619), .b(new_n14613), .O(new_n14942));
  inv1 g14749(.a(new_n14942), .O(new_n14943));
  nor2 g14750(.a(new_n14728), .b(new_n14722), .O(new_n14944));
  inv1 g14751(.a(new_n14944), .O(new_n14945));
  nor2 g14752(.a(new_n14673), .b(new_n14667), .O(new_n14946));
  inv1 g14753(.a(new_n14946), .O(new_n14947));
  nor2 g14754(.a(new_n14947), .b(new_n14945), .O(new_n14948));
  nor2 g14755(.a(new_n14946), .b(new_n14944), .O(new_n14949));
  nor2 g14756(.a(new_n14949), .b(new_n14948), .O(new_n14950));
  nor2 g14757(.a(new_n14849), .b(new_n14842), .O(new_n14951));
  inv1 g14758(.a(new_n14951), .O(new_n14952));
  nor2 g14759(.a(new_n14952), .b(new_n14950), .O(new_n14953));
  inv1 g14760(.a(new_n14950), .O(new_n14954));
  nor2 g14761(.a(new_n14951), .b(new_n14954), .O(new_n14955));
  nor2 g14762(.a(new_n14955), .b(new_n14953), .O(new_n14956));
  nor2 g14763(.a(new_n14781), .b(new_n14777), .O(new_n14957));
  inv1 g14764(.a(new_n14957), .O(new_n14958));
  nor2 g14765(.a(new_n14958), .b(new_n14956), .O(new_n14959));
  inv1 g14766(.a(new_n14956), .O(new_n14960));
  nor2 g14767(.a(new_n14957), .b(new_n14960), .O(new_n14961));
  nor2 g14768(.a(new_n14961), .b(new_n14959), .O(new_n14962));
  inv1 g14769(.a(new_n14962), .O(new_n14963));
  nor2 g14770(.a(new_n14772), .b(new_n14756), .O(new_n14964));
  nor2 g14771(.a(new_n10468), .b(new_n613), .O(new_n14965));
  inv1 g14772(.a(new_n14965), .O(new_n14966));
  nor2 g14773(.a(new_n14744), .b(new_n14737), .O(new_n14967));
  inv1 g14774(.a(new_n14967), .O(new_n14968));
  nor2 g14775(.a(new_n14968), .b(new_n14966), .O(new_n14969));
  nor2 g14776(.a(new_n14967), .b(new_n14965), .O(new_n14970));
  nor2 g14777(.a(new_n14970), .b(new_n14969), .O(new_n14971));
  nor2 g14778(.a(new_n14817), .b(new_n14810), .O(new_n14972));
  nor2 g14779(.a(new_n14972), .b(new_n14971), .O(new_n14973));
  inv1 g14780(.a(new_n14971), .O(new_n14974));
  inv1 g14781(.a(new_n14972), .O(new_n14975));
  nor2 g14782(.a(new_n14975), .b(new_n14974), .O(new_n14976));
  nor2 g14783(.a(new_n14976), .b(new_n14973), .O(new_n14977));
  inv1 g14784(.a(new_n14977), .O(new_n14978));
  nor2 g14785(.a(new_n14720), .b(new_n14713), .O(new_n14979));
  nor2 g14786(.a(new_n14704), .b(new_n14697), .O(new_n14980));
  nor2 g14787(.a(new_n14980), .b(new_n14979), .O(new_n14981));
  inv1 g14788(.a(new_n14979), .O(new_n14982));
  inv1 g14789(.a(new_n14980), .O(new_n14983));
  nor2 g14790(.a(new_n14983), .b(new_n14982), .O(new_n14984));
  nor2 g14791(.a(new_n14984), .b(new_n14981), .O(new_n14985));
  nor2 g14792(.a(new_n14770), .b(new_n14763), .O(new_n14986));
  nor2 g14793(.a(new_n14986), .b(new_n14985), .O(new_n14987));
  inv1 g14794(.a(new_n14985), .O(new_n14988));
  inv1 g14795(.a(new_n14986), .O(new_n14989));
  nor2 g14796(.a(new_n14989), .b(new_n14988), .O(new_n14990));
  nor2 g14797(.a(new_n14990), .b(new_n14987), .O(new_n14991));
  inv1 g14798(.a(new_n14991), .O(new_n14992));
  nor2 g14799(.a(new_n14992), .b(new_n14978), .O(new_n14993));
  nor2 g14800(.a(new_n14991), .b(new_n14977), .O(new_n14994));
  nor2 g14801(.a(new_n14994), .b(new_n14993), .O(new_n14995));
  inv1 g14802(.a(new_n14995), .O(new_n14996));
  nor2 g14803(.a(new_n14996), .b(new_n14964), .O(new_n14997));
  inv1 g14804(.a(new_n14964), .O(new_n14998));
  nor2 g14805(.a(new_n14995), .b(new_n14998), .O(new_n14999));
  nor2 g14806(.a(new_n14999), .b(new_n14997), .O(new_n15000));
  inv1 g14807(.a(new_n15000), .O(new_n15001));
  nor2 g14808(.a(new_n15001), .b(new_n14963), .O(new_n15002));
  nor2 g14809(.a(new_n15000), .b(new_n14962), .O(new_n15003));
  nor2 g14810(.a(new_n15003), .b(new_n15002), .O(new_n15004));
  nor2 g14811(.a(new_n15004), .b(new_n14943), .O(new_n15005));
  inv1 g14812(.a(new_n15004), .O(new_n15006));
  nor2 g14813(.a(new_n15006), .b(new_n14942), .O(new_n15007));
  nor2 g14814(.a(new_n15007), .b(new_n15005), .O(new_n15008));
  inv1 g14815(.a(new_n15008), .O(new_n15009));
  nor2 g14816(.a(new_n14640), .b(new_n14634), .O(new_n15010));
  inv1 g14817(.a(new_n15010), .O(new_n15011));
  nor2 g14818(.a(new_n8170), .b(new_n1297), .O(new_n15012));
  nor2 g14819(.a(new_n8026), .b(new_n1425), .O(new_n15013));
  nor2 g14820(.a(new_n15013), .b(new_n15012), .O(new_n15014));
  nor2 g14821(.a(new_n8170), .b(new_n1425), .O(new_n15015));
  inv1 g14822(.a(new_n15015), .O(new_n15016));
  nor2 g14823(.a(new_n15016), .b(new_n14395), .O(new_n15017));
  nor2 g14824(.a(new_n15017), .b(new_n15014), .O(new_n15018));
  nor2 g14825(.a(new_n15018), .b(new_n14739), .O(new_n15019));
  inv1 g14826(.a(new_n15018), .O(new_n15020));
  nor2 g14827(.a(new_n15020), .b(new_n14738), .O(new_n15021));
  nor2 g14828(.a(new_n15021), .b(new_n15019), .O(new_n15022));
  inv1 g14829(.a(new_n15022), .O(new_n15023));
  nor2 g14830(.a(new_n8946), .b(new_n1086), .O(new_n15024));
  inv1 g14831(.a(new_n15024), .O(new_n15025));
  nor2 g14832(.a(new_n8476), .b(new_n1199), .O(new_n15026));
  nor2 g14833(.a(new_n6958), .b(new_n1736), .O(new_n15027));
  nor2 g14834(.a(new_n15027), .b(new_n15026), .O(new_n15028));
  inv1 g14835(.a(new_n13276), .O(new_n15029));
  nor2 g14836(.a(new_n8476), .b(new_n1736), .O(new_n15030));
  inv1 g14837(.a(new_n15030), .O(new_n15031));
  nor2 g14838(.a(new_n15031), .b(new_n15029), .O(new_n15032));
  nor2 g14839(.a(new_n15032), .b(new_n15028), .O(new_n15033));
  nor2 g14840(.a(new_n15033), .b(new_n15025), .O(new_n15034));
  inv1 g14841(.a(new_n15033), .O(new_n15035));
  nor2 g14842(.a(new_n15035), .b(new_n15024), .O(new_n15036));
  nor2 g14843(.a(new_n15036), .b(new_n15034), .O(new_n15037));
  nor2 g14844(.a(new_n7294), .b(new_n1647), .O(new_n15038));
  inv1 g14845(.a(new_n15038), .O(new_n15039));
  nor2 g14846(.a(new_n14699), .b(\a[37] ), .O(new_n15040));
  nor2 g14847(.a(new_n5666), .b(new_n11186), .O(new_n15041));
  nor2 g14848(.a(new_n15041), .b(new_n15040), .O(new_n15042));
  nor2 g14849(.a(new_n15042), .b(new_n15039), .O(new_n15043));
  nor2 g14850(.a(new_n15040), .b(new_n15039), .O(new_n15044));
  nor2 g14851(.a(new_n15044), .b(new_n15041), .O(new_n15045));
  inv1 g14852(.a(new_n15045), .O(new_n15046));
  nor2 g14853(.a(new_n15046), .b(new_n15040), .O(new_n15047));
  nor2 g14854(.a(new_n15047), .b(new_n15043), .O(new_n15048));
  nor2 g14855(.a(new_n15048), .b(new_n15037), .O(new_n15049));
  inv1 g14856(.a(new_n15037), .O(new_n15050));
  inv1 g14857(.a(new_n15048), .O(new_n15051));
  nor2 g14858(.a(new_n15051), .b(new_n15050), .O(new_n15052));
  nor2 g14859(.a(new_n15052), .b(new_n15049), .O(new_n15053));
  nor2 g14860(.a(new_n15053), .b(new_n15023), .O(new_n15054));
  inv1 g14861(.a(new_n15053), .O(new_n15055));
  nor2 g14862(.a(new_n15055), .b(new_n15022), .O(new_n15056));
  nor2 g14863(.a(new_n15056), .b(new_n15054), .O(new_n15057));
  inv1 g14864(.a(new_n15057), .O(new_n15058));
  nor2 g14865(.a(new_n10320), .b(new_n699), .O(new_n15059));
  nor2 g14866(.a(new_n9658), .b(new_n847), .O(new_n15060));
  nor2 g14867(.a(new_n15060), .b(new_n14823), .O(new_n15061));
  inv1 g14868(.a(new_n14821), .O(new_n15062));
  nor2 g14869(.a(new_n9873), .b(new_n847), .O(new_n15063));
  inv1 g14870(.a(new_n15063), .O(new_n15064));
  nor2 g14871(.a(new_n15064), .b(new_n15062), .O(new_n15065));
  nor2 g14872(.a(new_n15065), .b(new_n15061), .O(new_n15066));
  inv1 g14873(.a(new_n15066), .O(new_n15067));
  nor2 g14874(.a(new_n15067), .b(new_n15059), .O(new_n15068));
  inv1 g14875(.a(new_n15059), .O(new_n15069));
  nor2 g14876(.a(new_n15066), .b(new_n15069), .O(new_n15070));
  nor2 g14877(.a(new_n15070), .b(new_n15068), .O(new_n15071));
  inv1 g14878(.a(new_n15071), .O(new_n15072));
  nor2 g14879(.a(new_n14752), .b(new_n14749), .O(new_n15073));
  nor2 g14880(.a(new_n9156), .b(new_n941), .O(new_n15074));
  inv1 g14881(.a(new_n15074), .O(new_n15075));
  nor2 g14882(.a(new_n6570), .b(new_n2121), .O(new_n15076));
  nor2 g14883(.a(new_n6274), .b(new_n2184), .O(new_n15077));
  nor2 g14884(.a(new_n15077), .b(new_n15076), .O(new_n15078));
  nor2 g14885(.a(new_n6570), .b(new_n2184), .O(new_n15079));
  inv1 g14886(.a(new_n15079), .O(new_n15080));
  nor2 g14887(.a(new_n15080), .b(new_n14479), .O(new_n15081));
  nor2 g14888(.a(new_n15081), .b(new_n15078), .O(new_n15082));
  nor2 g14889(.a(new_n15082), .b(new_n15075), .O(new_n15083));
  inv1 g14890(.a(new_n15082), .O(new_n15084));
  nor2 g14891(.a(new_n15084), .b(new_n15074), .O(new_n15085));
  nor2 g14892(.a(new_n15085), .b(new_n15083), .O(new_n15086));
  nor2 g14893(.a(new_n15086), .b(new_n15073), .O(new_n15087));
  inv1 g14894(.a(new_n15073), .O(new_n15088));
  inv1 g14895(.a(new_n15086), .O(new_n15089));
  nor2 g14896(.a(new_n15089), .b(new_n15088), .O(new_n15090));
  nor2 g14897(.a(new_n15090), .b(new_n15087), .O(new_n15091));
  nor2 g14898(.a(new_n15091), .b(new_n15072), .O(new_n15092));
  inv1 g14899(.a(new_n15091), .O(new_n15093));
  nor2 g14900(.a(new_n15093), .b(new_n15071), .O(new_n15094));
  nor2 g14901(.a(new_n15094), .b(new_n15092), .O(new_n15095));
  inv1 g14902(.a(new_n15095), .O(new_n15096));
  nor2 g14903(.a(new_n15096), .b(new_n15058), .O(new_n15097));
  nor2 g14904(.a(new_n15095), .b(new_n15057), .O(new_n15098));
  nor2 g14905(.a(new_n15098), .b(new_n15097), .O(new_n15099));
  nor2 g14906(.a(new_n15099), .b(new_n15011), .O(new_n15100));
  inv1 g14907(.a(new_n15099), .O(new_n15101));
  nor2 g14908(.a(new_n15101), .b(new_n15010), .O(new_n15102));
  nor2 g14909(.a(new_n15102), .b(new_n15100), .O(new_n15103));
  inv1 g14910(.a(new_n15103), .O(new_n15104));
  nor2 g14911(.a(new_n14609), .b(new_n14601), .O(new_n15105));
  nor2 g14912(.a(new_n14840), .b(new_n14833), .O(new_n15106));
  nor2 g14913(.a(new_n14828), .b(new_n14822), .O(new_n15107));
  nor2 g14914(.a(new_n15107), .b(new_n15106), .O(new_n15108));
  inv1 g14915(.a(new_n15106), .O(new_n15109));
  inv1 g14916(.a(new_n15107), .O(new_n15110));
  nor2 g14917(.a(new_n15110), .b(new_n15109), .O(new_n15111));
  nor2 g14918(.a(new_n15111), .b(new_n15108), .O(new_n15112));
  nor2 g14919(.a(new_n14588), .b(new_n14581), .O(new_n15113));
  nor2 g14920(.a(new_n15113), .b(new_n15112), .O(new_n15114));
  inv1 g14921(.a(new_n15112), .O(new_n15115));
  inv1 g14922(.a(new_n15113), .O(new_n15116));
  nor2 g14923(.a(new_n15116), .b(new_n15115), .O(new_n15117));
  nor2 g14924(.a(new_n15117), .b(new_n15114), .O(new_n15118));
  nor2 g14925(.a(new_n14598), .b(new_n14591), .O(new_n15119));
  inv1 g14926(.a(new_n15119), .O(new_n15120));
  nor2 g14927(.a(new_n15120), .b(new_n15118), .O(new_n15121));
  inv1 g14928(.a(new_n15118), .O(new_n15122));
  nor2 g14929(.a(new_n15119), .b(new_n15122), .O(new_n15123));
  nor2 g14930(.a(new_n15123), .b(new_n15121), .O(new_n15124));
  nor2 g14931(.a(new_n10895), .b(new_n569), .O(new_n15125));
  nor2 g14932(.a(new_n15125), .b(new_n14371), .O(new_n15126));
  nor2 g14933(.a(new_n11596), .b(new_n569), .O(new_n15127));
  inv1 g14934(.a(new_n15127), .O(new_n15128));
  nor2 g14935(.a(new_n15128), .b(new_n14698), .O(new_n15129));
  nor2 g14936(.a(new_n15129), .b(new_n15126), .O(new_n15130));
  inv1 g14937(.a(new_n15130), .O(new_n15131));
  nor2 g14938(.a(new_n15131), .b(new_n14714), .O(new_n15132));
  nor2 g14939(.a(new_n15130), .b(new_n14715), .O(new_n15133));
  nor2 g14940(.a(new_n15133), .b(new_n15132), .O(new_n15134));
  nor2 g14941(.a(new_n5796), .b(new_n2506), .O(new_n15135));
  nor2 g14942(.a(new_n5393), .b(new_n2660), .O(new_n15136));
  nor2 g14943(.a(new_n15136), .b(new_n15135), .O(new_n15137));
  nor2 g14944(.a(new_n5796), .b(new_n2660), .O(new_n15138));
  inv1 g14945(.a(new_n15138), .O(new_n15139));
  nor2 g14946(.a(new_n15139), .b(new_n14512), .O(new_n15140));
  nor2 g14947(.a(new_n15140), .b(new_n15137), .O(new_n15141));
  nor2 g14948(.a(new_n15141), .b(new_n14835), .O(new_n15142));
  inv1 g14949(.a(new_n15141), .O(new_n15143));
  nor2 g14950(.a(new_n15143), .b(new_n14834), .O(new_n15144));
  nor2 g14951(.a(new_n15144), .b(new_n15142), .O(new_n15145));
  nor2 g14952(.a(new_n15145), .b(new_n15134), .O(new_n15146));
  inv1 g14953(.a(new_n15134), .O(new_n15147));
  inv1 g14954(.a(new_n15145), .O(new_n15148));
  nor2 g14955(.a(new_n15148), .b(new_n15147), .O(new_n15149));
  nor2 g14956(.a(new_n15149), .b(new_n15146), .O(new_n15150));
  inv1 g14957(.a(new_n15150), .O(new_n15151));
  nor2 g14958(.a(new_n4366), .b(new_n3722), .O(new_n15152));
  nor2 g14959(.a(new_n4093), .b(new_n3870), .O(new_n15153));
  nor2 g14960(.a(new_n15153), .b(new_n15152), .O(new_n15154));
  nor2 g14961(.a(new_n4366), .b(new_n3870), .O(new_n15155));
  inv1 g14962(.a(new_n15155), .O(new_n15156));
  nor2 g14963(.a(new_n15156), .b(new_n14734), .O(new_n15157));
  nor2 g14964(.a(new_n15157), .b(new_n15154), .O(new_n15158));
  nor2 g14965(.a(new_n15158), .b(new_n14812), .O(new_n15159));
  inv1 g14966(.a(new_n15158), .O(new_n15160));
  nor2 g14967(.a(new_n15160), .b(new_n14811), .O(new_n15161));
  nor2 g14968(.a(new_n15161), .b(new_n15159), .O(new_n15162));
  nor2 g14969(.a(new_n15162), .b(new_n15151), .O(new_n15163));
  inv1 g14970(.a(new_n15162), .O(new_n15164));
  nor2 g14971(.a(new_n15164), .b(new_n15150), .O(new_n15165));
  nor2 g14972(.a(new_n15165), .b(new_n15163), .O(new_n15166));
  nor2 g14973(.a(new_n15166), .b(new_n15124), .O(new_n15167));
  inv1 g14974(.a(new_n15124), .O(new_n15168));
  inv1 g14975(.a(new_n15166), .O(new_n15169));
  nor2 g14976(.a(new_n15169), .b(new_n15168), .O(new_n15170));
  nor2 g14977(.a(new_n15170), .b(new_n15167), .O(new_n15171));
  inv1 g14978(.a(new_n15171), .O(new_n15172));
  nor2 g14979(.a(new_n15172), .b(new_n15105), .O(new_n15173));
  inv1 g14980(.a(new_n15105), .O(new_n15174));
  nor2 g14981(.a(new_n15171), .b(new_n15174), .O(new_n15175));
  nor2 g14982(.a(new_n15175), .b(new_n15173), .O(new_n15176));
  inv1 g14983(.a(new_n15176), .O(new_n15177));
  nor2 g14984(.a(new_n15177), .b(new_n15104), .O(new_n15178));
  nor2 g14985(.a(new_n15176), .b(new_n15103), .O(new_n15179));
  nor2 g14986(.a(new_n15179), .b(new_n15178), .O(new_n15180));
  inv1 g14987(.a(new_n15180), .O(new_n15181));
  nor2 g14988(.a(new_n15181), .b(new_n15009), .O(new_n15182));
  nor2 g14989(.a(new_n15180), .b(new_n15008), .O(new_n15183));
  nor2 g14990(.a(new_n15183), .b(new_n15182), .O(new_n15184));
  nor2 g14991(.a(new_n15184), .b(new_n14941), .O(new_n15185));
  inv1 g14992(.a(new_n14941), .O(new_n15186));
  inv1 g14993(.a(new_n15184), .O(new_n15187));
  nor2 g14994(.a(new_n15187), .b(new_n15186), .O(new_n15188));
  nor2 g14995(.a(new_n15188), .b(new_n15185), .O(new_n15189));
  nor2 g14996(.a(new_n15189), .b(new_n14888), .O(new_n15190));
  inv1 g14997(.a(new_n15189), .O(new_n15191));
  nor2 g14998(.a(new_n15191), .b(new_n14887), .O(new_n15192));
  nor2 g14999(.a(new_n15192), .b(new_n15190), .O(new_n15193));
  inv1 g15000(.a(new_n15193), .O(new_n15194));
  nor2 g15001(.a(new_n14884), .b(new_n14876), .O(new_n15195));
  nor2 g15002(.a(new_n15195), .b(new_n15194), .O(new_n15196));
  inv1 g15003(.a(new_n15195), .O(new_n15197));
  nor2 g15004(.a(new_n15197), .b(new_n15193), .O(new_n15198));
  nor2 g15005(.a(new_n15198), .b(new_n15196), .O(new_n15199));
  inv1 g15006(.a(new_n15199), .O(\asquared[74] ));
  nor2 g15007(.a(new_n15188), .b(new_n14940), .O(new_n15201));
  inv1 g15008(.a(new_n15201), .O(new_n15202));
  nor2 g15009(.a(new_n15182), .b(new_n15007), .O(new_n15203));
  nor2 g15010(.a(new_n15178), .b(new_n15173), .O(new_n15204));
  nor2 g15011(.a(new_n15002), .b(new_n14961), .O(new_n15205));
  nor2 g15012(.a(new_n14990), .b(new_n14984), .O(new_n15206));
  inv1 g15013(.a(new_n15206), .O(new_n15207));
  nor2 g15014(.a(new_n14976), .b(new_n14969), .O(new_n15208));
  inv1 g15015(.a(new_n15208), .O(new_n15209));
  nor2 g15016(.a(new_n15209), .b(new_n15207), .O(new_n15210));
  nor2 g15017(.a(new_n15208), .b(new_n15206), .O(new_n15211));
  nor2 g15018(.a(new_n15211), .b(new_n15210), .O(new_n15212));
  nor2 g15019(.a(new_n15094), .b(new_n15087), .O(new_n15213));
  inv1 g15020(.a(new_n15213), .O(new_n15214));
  nor2 g15021(.a(new_n15214), .b(new_n15212), .O(new_n15215));
  inv1 g15022(.a(new_n15212), .O(new_n15216));
  nor2 g15023(.a(new_n15213), .b(new_n15216), .O(new_n15217));
  nor2 g15024(.a(new_n15217), .b(new_n15215), .O(new_n15218));
  inv1 g15025(.a(new_n15218), .O(new_n15219));
  nor2 g15026(.a(new_n14997), .b(new_n14993), .O(new_n15220));
  inv1 g15027(.a(new_n15220), .O(new_n15221));
  nor2 g15028(.a(new_n14955), .b(new_n14949), .O(new_n15222));
  inv1 g15029(.a(new_n15222), .O(new_n15223));
  nor2 g15030(.a(new_n15223), .b(new_n15221), .O(new_n15224));
  nor2 g15031(.a(new_n15222), .b(new_n15220), .O(new_n15225));
  nor2 g15032(.a(new_n15225), .b(new_n15224), .O(new_n15226));
  inv1 g15033(.a(new_n15226), .O(new_n15227));
  nor2 g15034(.a(new_n15227), .b(new_n15219), .O(new_n15228));
  nor2 g15035(.a(new_n15226), .b(new_n15218), .O(new_n15229));
  nor2 g15036(.a(new_n15229), .b(new_n15228), .O(new_n15230));
  inv1 g15037(.a(new_n15230), .O(new_n15231));
  nor2 g15038(.a(new_n15231), .b(new_n15205), .O(new_n15232));
  inv1 g15039(.a(new_n15205), .O(new_n15233));
  nor2 g15040(.a(new_n15230), .b(new_n15233), .O(new_n15234));
  nor2 g15041(.a(new_n15234), .b(new_n15232), .O(new_n15235));
  inv1 g15042(.a(new_n15235), .O(new_n15236));
  nor2 g15043(.a(new_n15236), .b(new_n15204), .O(new_n15237));
  inv1 g15044(.a(new_n15204), .O(new_n15238));
  nor2 g15045(.a(new_n15235), .b(new_n15238), .O(new_n15239));
  nor2 g15046(.a(new_n15239), .b(new_n15237), .O(new_n15240));
  inv1 g15047(.a(new_n15240), .O(new_n15241));
  nor2 g15048(.a(new_n15241), .b(new_n15203), .O(new_n15242));
  inv1 g15049(.a(new_n15203), .O(new_n15243));
  nor2 g15050(.a(new_n15240), .b(new_n15243), .O(new_n15244));
  nor2 g15051(.a(new_n15244), .b(new_n15242), .O(new_n15245));
  inv1 g15052(.a(new_n15245), .O(new_n15246));
  nor2 g15053(.a(new_n14934), .b(new_n14929), .O(new_n15247));
  nor2 g15054(.a(new_n15161), .b(new_n15154), .O(new_n15248));
  nor2 g15055(.a(new_n14906), .b(new_n14899), .O(new_n15249));
  nor2 g15056(.a(new_n15249), .b(new_n15248), .O(new_n15250));
  inv1 g15057(.a(new_n15248), .O(new_n15251));
  inv1 g15058(.a(new_n15249), .O(new_n15252));
  nor2 g15059(.a(new_n15252), .b(new_n15251), .O(new_n15253));
  nor2 g15060(.a(new_n15253), .b(new_n15250), .O(new_n15254));
  inv1 g15061(.a(new_n15254), .O(new_n15255));
  nor2 g15062(.a(new_n10468), .b(new_n699), .O(new_n15256));
  inv1 g15063(.a(new_n15256), .O(new_n15257));
  nor2 g15064(.a(new_n10320), .b(new_n800), .O(new_n15258));
  nor2 g15065(.a(new_n15258), .b(new_n15063), .O(new_n15259));
  nor2 g15066(.a(new_n10320), .b(new_n847), .O(new_n15260));
  inv1 g15067(.a(new_n15260), .O(new_n15261));
  nor2 g15068(.a(new_n15261), .b(new_n14824), .O(new_n15262));
  nor2 g15069(.a(new_n15262), .b(new_n15259), .O(new_n15263));
  nor2 g15070(.a(new_n15263), .b(new_n15257), .O(new_n15264));
  inv1 g15071(.a(new_n15263), .O(new_n15265));
  nor2 g15072(.a(new_n15265), .b(new_n15256), .O(new_n15266));
  nor2 g15073(.a(new_n15266), .b(new_n15264), .O(new_n15267));
  nor2 g15074(.a(new_n15267), .b(new_n15255), .O(new_n15268));
  inv1 g15075(.a(new_n15267), .O(new_n15269));
  nor2 g15076(.a(new_n15269), .b(new_n15254), .O(new_n15270));
  nor2 g15077(.a(new_n15270), .b(new_n15268), .O(new_n15271));
  nor2 g15078(.a(new_n15056), .b(new_n15049), .O(new_n15272));
  inv1 g15079(.a(new_n15272), .O(new_n15273));
  nor2 g15080(.a(new_n15273), .b(new_n15271), .O(new_n15274));
  inv1 g15081(.a(new_n15271), .O(new_n15275));
  nor2 g15082(.a(new_n15272), .b(new_n15275), .O(new_n15276));
  nor2 g15083(.a(new_n15276), .b(new_n15274), .O(new_n15277));
  nor2 g15084(.a(new_n14915), .b(new_n14908), .O(new_n15278));
  inv1 g15085(.a(new_n15278), .O(new_n15279));
  nor2 g15086(.a(new_n15279), .b(new_n15277), .O(new_n15280));
  inv1 g15087(.a(new_n15277), .O(new_n15281));
  nor2 g15088(.a(new_n15278), .b(new_n15281), .O(new_n15282));
  nor2 g15089(.a(new_n15282), .b(new_n15280), .O(new_n15283));
  inv1 g15090(.a(new_n15283), .O(new_n15284));
  nor2 g15091(.a(new_n15102), .b(new_n15097), .O(new_n15285));
  nor2 g15092(.a(new_n15170), .b(new_n15123), .O(new_n15286));
  nor2 g15093(.a(new_n15286), .b(new_n15285), .O(new_n15287));
  inv1 g15094(.a(new_n15285), .O(new_n15288));
  inv1 g15095(.a(new_n15286), .O(new_n15289));
  nor2 g15096(.a(new_n15289), .b(new_n15288), .O(new_n15290));
  nor2 g15097(.a(new_n15290), .b(new_n15287), .O(new_n15291));
  inv1 g15098(.a(new_n15291), .O(new_n15292));
  nor2 g15099(.a(new_n15292), .b(new_n15284), .O(new_n15293));
  nor2 g15100(.a(new_n15291), .b(new_n15283), .O(new_n15294));
  nor2 g15101(.a(new_n15294), .b(new_n15293), .O(new_n15295));
  inv1 g15102(.a(new_n15295), .O(new_n15296));
  nor2 g15103(.a(new_n15296), .b(new_n15247), .O(new_n15297));
  inv1 g15104(.a(new_n15247), .O(new_n15298));
  nor2 g15105(.a(new_n15295), .b(new_n15298), .O(new_n15299));
  nor2 g15106(.a(new_n15299), .b(new_n15297), .O(new_n15300));
  inv1 g15107(.a(new_n15300), .O(new_n15301));
  nor2 g15108(.a(new_n14924), .b(new_n14919), .O(new_n15302));
  nor2 g15109(.a(new_n15085), .b(new_n15078), .O(new_n15303));
  nor2 g15110(.a(new_n15144), .b(new_n15137), .O(new_n15304));
  nor2 g15111(.a(new_n15304), .b(new_n15303), .O(new_n15305));
  inv1 g15112(.a(new_n15303), .O(new_n15306));
  inv1 g15113(.a(new_n15304), .O(new_n15307));
  nor2 g15114(.a(new_n15307), .b(new_n15306), .O(new_n15308));
  nor2 g15115(.a(new_n15308), .b(new_n15305), .O(new_n15309));
  nor2 g15116(.a(new_n15068), .b(new_n15061), .O(new_n15310));
  nor2 g15117(.a(new_n15310), .b(new_n15309), .O(new_n15311));
  inv1 g15118(.a(new_n15309), .O(new_n15312));
  inv1 g15119(.a(new_n15310), .O(new_n15313));
  nor2 g15120(.a(new_n15313), .b(new_n15312), .O(new_n15314));
  nor2 g15121(.a(new_n15314), .b(new_n15311), .O(new_n15315));
  inv1 g15122(.a(new_n15315), .O(new_n15316));
  nor2 g15123(.a(new_n15036), .b(new_n15028), .O(new_n15317));
  nor2 g15124(.a(new_n15021), .b(new_n15014), .O(new_n15318));
  nor2 g15125(.a(new_n15318), .b(new_n15317), .O(new_n15319));
  inv1 g15126(.a(new_n15317), .O(new_n15320));
  inv1 g15127(.a(new_n15318), .O(new_n15321));
  nor2 g15128(.a(new_n15321), .b(new_n15320), .O(new_n15322));
  nor2 g15129(.a(new_n15322), .b(new_n15319), .O(new_n15323));
  nor2 g15130(.a(new_n15132), .b(new_n15126), .O(new_n15324));
  nor2 g15131(.a(new_n15324), .b(new_n15323), .O(new_n15325));
  inv1 g15132(.a(new_n15323), .O(new_n15326));
  inv1 g15133(.a(new_n15324), .O(new_n15327));
  nor2 g15134(.a(new_n15327), .b(new_n15326), .O(new_n15328));
  nor2 g15135(.a(new_n15328), .b(new_n15325), .O(new_n15329));
  nor2 g15136(.a(new_n15163), .b(new_n15146), .O(new_n15330));
  inv1 g15137(.a(new_n15330), .O(new_n15331));
  nor2 g15138(.a(new_n15331), .b(new_n15329), .O(new_n15332));
  inv1 g15139(.a(new_n15329), .O(new_n15333));
  nor2 g15140(.a(new_n15330), .b(new_n15333), .O(new_n15334));
  nor2 g15141(.a(new_n15334), .b(new_n15332), .O(new_n15335));
  inv1 g15142(.a(new_n15335), .O(new_n15336));
  nor2 g15143(.a(new_n15336), .b(new_n15316), .O(new_n15337));
  nor2 g15144(.a(new_n15335), .b(new_n15315), .O(new_n15338));
  nor2 g15145(.a(new_n15338), .b(new_n15337), .O(new_n15339));
  inv1 g15146(.a(new_n15339), .O(new_n15340));
  nor2 g15147(.a(new_n15340), .b(new_n15302), .O(new_n15341));
  inv1 g15148(.a(new_n15302), .O(new_n15342));
  nor2 g15149(.a(new_n15339), .b(new_n15342), .O(new_n15343));
  nor2 g15150(.a(new_n15343), .b(new_n15341), .O(new_n15344));
  inv1 g15151(.a(new_n15344), .O(new_n15345));
  nor2 g15152(.a(new_n15117), .b(new_n15111), .O(new_n15346));
  inv1 g15153(.a(new_n15346), .O(new_n15347));
  nor2 g15154(.a(new_n5971), .b(new_n2506), .O(new_n15348));
  inv1 g15155(.a(new_n15348), .O(new_n15349));
  nor2 g15156(.a(new_n15138), .b(new_n12032), .O(new_n15350));
  nor2 g15157(.a(new_n15139), .b(new_n12033), .O(new_n15351));
  nor2 g15158(.a(new_n15351), .b(new_n15350), .O(new_n15352));
  nor2 g15159(.a(new_n15352), .b(new_n15349), .O(new_n15353));
  inv1 g15160(.a(new_n15352), .O(new_n15354));
  nor2 g15161(.a(new_n15354), .b(new_n15348), .O(new_n15355));
  nor2 g15162(.a(new_n15355), .b(new_n15353), .O(new_n15356));
  nor2 g15163(.a(new_n10895), .b(new_n613), .O(new_n15357));
  nor2 g15164(.a(new_n11186), .b(new_n569), .O(new_n15358));
  nor2 g15165(.a(new_n15358), .b(new_n15357), .O(new_n15359));
  inv1 g15166(.a(new_n15125), .O(new_n15360));
  nor2 g15167(.a(new_n11186), .b(new_n613), .O(new_n15361));
  inv1 g15168(.a(new_n15361), .O(new_n15362));
  nor2 g15169(.a(new_n15362), .b(new_n15360), .O(new_n15363));
  nor2 g15170(.a(new_n15363), .b(new_n15359), .O(new_n15364));
  inv1 g15171(.a(new_n15364), .O(new_n15365));
  nor2 g15172(.a(new_n15365), .b(new_n15045), .O(new_n15366));
  nor2 g15173(.a(new_n15364), .b(new_n15046), .O(new_n15367));
  nor2 g15174(.a(new_n15367), .b(new_n15366), .O(new_n15368));
  inv1 g15175(.a(new_n15368), .O(new_n15369));
  nor2 g15176(.a(new_n15369), .b(new_n15356), .O(new_n15370));
  inv1 g15177(.a(new_n15356), .O(new_n15371));
  nor2 g15178(.a(new_n15368), .b(new_n15371), .O(new_n15372));
  nor2 g15179(.a(new_n15372), .b(new_n15370), .O(new_n15373));
  nor2 g15180(.a(new_n15373), .b(new_n15347), .O(new_n15374));
  inv1 g15181(.a(new_n15373), .O(new_n15375));
  nor2 g15182(.a(new_n15375), .b(new_n15346), .O(new_n15376));
  nor2 g15183(.a(new_n15376), .b(new_n15374), .O(new_n15377));
  inv1 g15184(.a(new_n15377), .O(new_n15378));
  nor2 g15185(.a(new_n6893), .b(new_n2121), .O(new_n15379));
  inv1 g15186(.a(new_n15379), .O(new_n15380));
  nor2 g15187(.a(new_n6274), .b(new_n2433), .O(new_n15381));
  nor2 g15188(.a(new_n15381), .b(new_n15079), .O(new_n15382));
  inv1 g15189(.a(new_n15077), .O(new_n15383));
  nor2 g15190(.a(new_n6570), .b(new_n2433), .O(new_n15384));
  inv1 g15191(.a(new_n15384), .O(new_n15385));
  nor2 g15192(.a(new_n15385), .b(new_n15383), .O(new_n15386));
  nor2 g15193(.a(new_n15386), .b(new_n15382), .O(new_n15387));
  nor2 g15194(.a(new_n15387), .b(new_n15380), .O(new_n15388));
  inv1 g15195(.a(new_n15387), .O(new_n15389));
  nor2 g15196(.a(new_n15389), .b(new_n15379), .O(new_n15390));
  nor2 g15197(.a(new_n15390), .b(new_n15388), .O(new_n15391));
  inv1 g15198(.a(new_n15391), .O(new_n15392));
  nor2 g15199(.a(new_n11596), .b(new_n502), .O(new_n15393));
  nor2 g15200(.a(new_n5393), .b(new_n2826), .O(new_n15394));
  nor2 g15201(.a(new_n5178), .b(new_n3057), .O(new_n15395));
  nor2 g15202(.a(new_n15395), .b(new_n15394), .O(new_n15396));
  nor2 g15203(.a(new_n5393), .b(new_n3057), .O(new_n15397));
  inv1 g15204(.a(new_n15397), .O(new_n15398));
  nor2 g15205(.a(new_n15398), .b(new_n14583), .O(new_n15399));
  nor2 g15206(.a(new_n15399), .b(new_n15396), .O(new_n15400));
  inv1 g15207(.a(new_n15400), .O(new_n15401));
  nor2 g15208(.a(new_n15401), .b(new_n15393), .O(new_n15402));
  inv1 g15209(.a(new_n15393), .O(new_n15403));
  nor2 g15210(.a(new_n15400), .b(new_n15403), .O(new_n15404));
  nor2 g15211(.a(new_n15404), .b(new_n15402), .O(new_n15405));
  nor2 g15212(.a(new_n9156), .b(new_n1086), .O(new_n15406));
  nor2 g15213(.a(new_n6958), .b(new_n1903), .O(new_n15407));
  nor2 g15214(.a(new_n15407), .b(new_n15406), .O(new_n15408));
  nor2 g15215(.a(new_n9156), .b(new_n1903), .O(new_n15409));
  inv1 g15216(.a(new_n15409), .O(new_n15410));
  nor2 g15217(.a(new_n15410), .b(new_n13126), .O(new_n15411));
  nor2 g15218(.a(new_n15411), .b(new_n15408), .O(new_n15412));
  nor2 g15219(.a(new_n15412), .b(new_n14901), .O(new_n15413));
  inv1 g15220(.a(new_n15412), .O(new_n15414));
  nor2 g15221(.a(new_n15414), .b(new_n14900), .O(new_n15415));
  nor2 g15222(.a(new_n15415), .b(new_n15413), .O(new_n15416));
  nor2 g15223(.a(new_n15416), .b(new_n15405), .O(new_n15417));
  inv1 g15224(.a(new_n15405), .O(new_n15418));
  inv1 g15225(.a(new_n15416), .O(new_n15419));
  nor2 g15226(.a(new_n15419), .b(new_n15418), .O(new_n15420));
  nor2 g15227(.a(new_n15420), .b(new_n15417), .O(new_n15421));
  nor2 g15228(.a(new_n15421), .b(new_n15392), .O(new_n15422));
  inv1 g15229(.a(new_n15421), .O(new_n15423));
  nor2 g15230(.a(new_n15423), .b(new_n15391), .O(new_n15424));
  nor2 g15231(.a(new_n15424), .b(new_n15422), .O(new_n15425));
  inv1 g15232(.a(new_n15425), .O(new_n15426));
  nor2 g15233(.a(new_n7537), .b(new_n1647), .O(new_n15427));
  nor2 g15234(.a(new_n7294), .b(new_n1736), .O(new_n15428));
  nor2 g15235(.a(new_n15428), .b(new_n15427), .O(new_n15429));
  nor2 g15236(.a(new_n7537), .b(new_n1736), .O(new_n15430));
  inv1 g15237(.a(new_n15430), .O(new_n15431));
  nor2 g15238(.a(new_n15431), .b(new_n15039), .O(new_n15432));
  nor2 g15239(.a(new_n15432), .b(new_n15429), .O(new_n15433));
  nor2 g15240(.a(new_n15433), .b(new_n15156), .O(new_n15434));
  inv1 g15241(.a(new_n15433), .O(new_n15435));
  nor2 g15242(.a(new_n15435), .b(new_n15155), .O(new_n15436));
  nor2 g15243(.a(new_n15436), .b(new_n15434), .O(new_n15437));
  inv1 g15244(.a(new_n15437), .O(new_n15438));
  nor2 g15245(.a(new_n8026), .b(new_n1493), .O(new_n15439));
  nor2 g15246(.a(new_n15015), .b(new_n11747), .O(new_n15440));
  nor2 g15247(.a(new_n8946), .b(new_n1425), .O(new_n15441));
  inv1 g15248(.a(new_n15441), .O(new_n15442));
  nor2 g15249(.a(new_n15442), .b(new_n14807), .O(new_n15443));
  nor2 g15250(.a(new_n15443), .b(new_n15440), .O(new_n15444));
  inv1 g15251(.a(new_n15444), .O(new_n15445));
  nor2 g15252(.a(new_n15445), .b(new_n15439), .O(new_n15446));
  inv1 g15253(.a(new_n15439), .O(new_n15447));
  nor2 g15254(.a(new_n15444), .b(new_n15447), .O(new_n15448));
  nor2 g15255(.a(new_n15448), .b(new_n15446), .O(new_n15449));
  nor2 g15256(.a(new_n4425), .b(new_n3722), .O(new_n15450));
  nor2 g15257(.a(new_n4682), .b(new_n3533), .O(new_n15451));
  nor2 g15258(.a(new_n15451), .b(new_n15450), .O(new_n15452));
  nor2 g15259(.a(new_n4682), .b(new_n3722), .O(new_n15453));
  inv1 g15260(.a(new_n15453), .O(new_n15454));
  nor2 g15261(.a(new_n15454), .b(new_n14812), .O(new_n15455));
  nor2 g15262(.a(new_n15455), .b(new_n15452), .O(new_n15456));
  nor2 g15263(.a(new_n15456), .b(new_n14765), .O(new_n15457));
  inv1 g15264(.a(new_n15456), .O(new_n15458));
  nor2 g15265(.a(new_n15458), .b(new_n14764), .O(new_n15459));
  nor2 g15266(.a(new_n15459), .b(new_n15457), .O(new_n15460));
  nor2 g15267(.a(new_n15460), .b(new_n15449), .O(new_n15461));
  inv1 g15268(.a(new_n15449), .O(new_n15462));
  inv1 g15269(.a(new_n15460), .O(new_n15463));
  nor2 g15270(.a(new_n15463), .b(new_n15462), .O(new_n15464));
  nor2 g15271(.a(new_n15464), .b(new_n15461), .O(new_n15465));
  nor2 g15272(.a(new_n15465), .b(new_n15438), .O(new_n15466));
  inv1 g15273(.a(new_n15465), .O(new_n15467));
  nor2 g15274(.a(new_n15467), .b(new_n15437), .O(new_n15468));
  nor2 g15275(.a(new_n15468), .b(new_n15466), .O(new_n15469));
  inv1 g15276(.a(new_n15469), .O(new_n15470));
  nor2 g15277(.a(new_n15470), .b(new_n15426), .O(new_n15471));
  nor2 g15278(.a(new_n15469), .b(new_n15425), .O(new_n15472));
  nor2 g15279(.a(new_n15472), .b(new_n15471), .O(new_n15473));
  inv1 g15280(.a(new_n15473), .O(new_n15474));
  nor2 g15281(.a(new_n15474), .b(new_n15378), .O(new_n15475));
  nor2 g15282(.a(new_n15473), .b(new_n15377), .O(new_n15476));
  nor2 g15283(.a(new_n15476), .b(new_n15475), .O(new_n15477));
  inv1 g15284(.a(new_n15477), .O(new_n15478));
  nor2 g15285(.a(new_n15478), .b(new_n15345), .O(new_n15479));
  nor2 g15286(.a(new_n15477), .b(new_n15344), .O(new_n15480));
  nor2 g15287(.a(new_n15480), .b(new_n15479), .O(new_n15481));
  inv1 g15288(.a(new_n15481), .O(new_n15482));
  nor2 g15289(.a(new_n15482), .b(new_n15301), .O(new_n15483));
  nor2 g15290(.a(new_n15481), .b(new_n15300), .O(new_n15484));
  nor2 g15291(.a(new_n15484), .b(new_n15483), .O(new_n15485));
  inv1 g15292(.a(new_n15485), .O(new_n15486));
  nor2 g15293(.a(new_n15486), .b(new_n15246), .O(new_n15487));
  nor2 g15294(.a(new_n15485), .b(new_n15245), .O(new_n15488));
  nor2 g15295(.a(new_n15488), .b(new_n15487), .O(new_n15489));
  nor2 g15296(.a(new_n15489), .b(new_n15202), .O(new_n15490));
  inv1 g15297(.a(new_n15489), .O(new_n15491));
  nor2 g15298(.a(new_n15491), .b(new_n15201), .O(new_n15492));
  nor2 g15299(.a(new_n15492), .b(new_n15490), .O(new_n15493));
  nor2 g15300(.a(new_n15196), .b(new_n15190), .O(new_n15494));
  inv1 g15301(.a(new_n15494), .O(new_n15495));
  nor2 g15302(.a(new_n15495), .b(new_n15493), .O(new_n15496));
  inv1 g15303(.a(new_n15493), .O(new_n15497));
  nor2 g15304(.a(new_n15494), .b(new_n15497), .O(new_n15498));
  nor2 g15305(.a(new_n15498), .b(new_n15496), .O(new_n15499));
  inv1 g15306(.a(new_n15499), .O(\asquared[75] ));
  nor2 g15307(.a(new_n15487), .b(new_n15242), .O(new_n15501));
  nor2 g15308(.a(new_n15237), .b(new_n15232), .O(new_n15502));
  inv1 g15309(.a(new_n15502), .O(new_n15503));
  nor2 g15310(.a(new_n15328), .b(new_n15322), .O(new_n15504));
  inv1 g15311(.a(new_n15504), .O(new_n15505));
  nor2 g15312(.a(new_n15268), .b(new_n15253), .O(new_n15506));
  inv1 g15313(.a(new_n15506), .O(new_n15507));
  nor2 g15314(.a(new_n15507), .b(new_n15505), .O(new_n15508));
  nor2 g15315(.a(new_n15506), .b(new_n15504), .O(new_n15509));
  nor2 g15316(.a(new_n15509), .b(new_n15508), .O(new_n15510));
  nor2 g15317(.a(new_n15314), .b(new_n15308), .O(new_n15511));
  inv1 g15318(.a(new_n15511), .O(new_n15512));
  nor2 g15319(.a(new_n15512), .b(new_n15510), .O(new_n15513));
  inv1 g15320(.a(new_n15510), .O(new_n15514));
  nor2 g15321(.a(new_n15511), .b(new_n15514), .O(new_n15515));
  nor2 g15322(.a(new_n15515), .b(new_n15513), .O(new_n15516));
  inv1 g15323(.a(new_n15516), .O(new_n15517));
  nor2 g15324(.a(new_n15475), .b(new_n15471), .O(new_n15518));
  nor2 g15325(.a(new_n15518), .b(new_n15517), .O(new_n15519));
  inv1 g15326(.a(new_n15518), .O(new_n15520));
  nor2 g15327(.a(new_n15520), .b(new_n15516), .O(new_n15521));
  nor2 g15328(.a(new_n15521), .b(new_n15519), .O(new_n15522));
  inv1 g15329(.a(new_n15522), .O(new_n15523));
  nor2 g15330(.a(new_n15376), .b(new_n15370), .O(new_n15524));
  nor2 g15331(.a(new_n15459), .b(new_n15452), .O(new_n15525));
  nor2 g15332(.a(new_n15436), .b(new_n15429), .O(new_n15526));
  nor2 g15333(.a(new_n15526), .b(new_n15525), .O(new_n15527));
  inv1 g15334(.a(new_n15525), .O(new_n15528));
  inv1 g15335(.a(new_n15526), .O(new_n15529));
  nor2 g15336(.a(new_n15529), .b(new_n15528), .O(new_n15530));
  nor2 g15337(.a(new_n15530), .b(new_n15527), .O(new_n15531));
  nor2 g15338(.a(new_n15446), .b(new_n15440), .O(new_n15532));
  nor2 g15339(.a(new_n15532), .b(new_n15531), .O(new_n15533));
  inv1 g15340(.a(new_n15531), .O(new_n15534));
  inv1 g15341(.a(new_n15532), .O(new_n15535));
  nor2 g15342(.a(new_n15535), .b(new_n15534), .O(new_n15536));
  nor2 g15343(.a(new_n15536), .b(new_n15533), .O(new_n15537));
  inv1 g15344(.a(new_n15537), .O(new_n15538));
  nor2 g15345(.a(new_n15415), .b(new_n15408), .O(new_n15539));
  nor2 g15346(.a(new_n15402), .b(new_n15396), .O(new_n15540));
  nor2 g15347(.a(new_n15540), .b(new_n15539), .O(new_n15541));
  inv1 g15348(.a(new_n15539), .O(new_n15542));
  inv1 g15349(.a(new_n15540), .O(new_n15543));
  nor2 g15350(.a(new_n15543), .b(new_n15542), .O(new_n15544));
  nor2 g15351(.a(new_n15544), .b(new_n15541), .O(new_n15545));
  nor2 g15352(.a(new_n15366), .b(new_n15363), .O(new_n15546));
  inv1 g15353(.a(new_n15546), .O(new_n15547));
  nor2 g15354(.a(new_n15547), .b(new_n15545), .O(new_n15548));
  inv1 g15355(.a(new_n15545), .O(new_n15549));
  nor2 g15356(.a(new_n15546), .b(new_n15549), .O(new_n15550));
  nor2 g15357(.a(new_n15550), .b(new_n15548), .O(new_n15551));
  inv1 g15358(.a(new_n15551), .O(new_n15552));
  nor2 g15359(.a(new_n15552), .b(new_n15538), .O(new_n15553));
  nor2 g15360(.a(new_n15551), .b(new_n15537), .O(new_n15554));
  nor2 g15361(.a(new_n15554), .b(new_n15553), .O(new_n15555));
  inv1 g15362(.a(new_n15555), .O(new_n15556));
  nor2 g15363(.a(new_n15556), .b(new_n15524), .O(new_n15557));
  inv1 g15364(.a(new_n15524), .O(new_n15558));
  nor2 g15365(.a(new_n15555), .b(new_n15558), .O(new_n15559));
  nor2 g15366(.a(new_n15559), .b(new_n15557), .O(new_n15560));
  inv1 g15367(.a(new_n15560), .O(new_n15561));
  nor2 g15368(.a(new_n15561), .b(new_n15523), .O(new_n15562));
  nor2 g15369(.a(new_n15560), .b(new_n15522), .O(new_n15563));
  nor2 g15370(.a(new_n15563), .b(new_n15562), .O(new_n15564));
  nor2 g15371(.a(new_n15564), .b(new_n15503), .O(new_n15565));
  inv1 g15372(.a(new_n15564), .O(new_n15566));
  nor2 g15373(.a(new_n15566), .b(new_n15502), .O(new_n15567));
  nor2 g15374(.a(new_n15567), .b(new_n15565), .O(new_n15568));
  nor2 g15375(.a(new_n15228), .b(new_n15225), .O(new_n15569));
  nor2 g15376(.a(new_n15355), .b(new_n15350), .O(new_n15570));
  nor2 g15377(.a(new_n15390), .b(new_n15382), .O(new_n15571));
  nor2 g15378(.a(new_n15571), .b(new_n15570), .O(new_n15572));
  inv1 g15379(.a(new_n15570), .O(new_n15573));
  inv1 g15380(.a(new_n15571), .O(new_n15574));
  nor2 g15381(.a(new_n15574), .b(new_n15573), .O(new_n15575));
  nor2 g15382(.a(new_n15575), .b(new_n15572), .O(new_n15576));
  nor2 g15383(.a(new_n15266), .b(new_n15259), .O(new_n15577));
  nor2 g15384(.a(new_n15577), .b(new_n15576), .O(new_n15578));
  inv1 g15385(.a(new_n15576), .O(new_n15579));
  inv1 g15386(.a(new_n15577), .O(new_n15580));
  nor2 g15387(.a(new_n15580), .b(new_n15579), .O(new_n15581));
  nor2 g15388(.a(new_n15581), .b(new_n15578), .O(new_n15582));
  inv1 g15389(.a(new_n15582), .O(new_n15583));
  nor2 g15390(.a(new_n15468), .b(new_n15461), .O(new_n15584));
  inv1 g15391(.a(new_n15584), .O(new_n15585));
  nor2 g15392(.a(new_n15424), .b(new_n15417), .O(new_n15586));
  inv1 g15393(.a(new_n15586), .O(new_n15587));
  nor2 g15394(.a(new_n15587), .b(new_n15585), .O(new_n15588));
  nor2 g15395(.a(new_n15586), .b(new_n15584), .O(new_n15589));
  nor2 g15396(.a(new_n15589), .b(new_n15588), .O(new_n15590));
  inv1 g15397(.a(new_n15590), .O(new_n15591));
  nor2 g15398(.a(new_n15591), .b(new_n15583), .O(new_n15592));
  nor2 g15399(.a(new_n15590), .b(new_n15582), .O(new_n15593));
  nor2 g15400(.a(new_n15593), .b(new_n15592), .O(new_n15594));
  inv1 g15401(.a(new_n15594), .O(new_n15595));
  nor2 g15402(.a(new_n15595), .b(new_n15569), .O(new_n15596));
  inv1 g15403(.a(new_n15569), .O(new_n15597));
  nor2 g15404(.a(new_n15594), .b(new_n15597), .O(new_n15598));
  nor2 g15405(.a(new_n15598), .b(new_n15596), .O(new_n15599));
  inv1 g15406(.a(new_n15599), .O(new_n15600));
  nor2 g15407(.a(new_n15217), .b(new_n15211), .O(new_n15601));
  inv1 g15408(.a(new_n15601), .O(new_n15602));
  nor2 g15409(.a(new_n5971), .b(new_n2660), .O(new_n15603));
  nor2 g15410(.a(new_n9156), .b(new_n1199), .O(new_n15604));
  nor2 g15411(.a(new_n15604), .b(new_n15127), .O(new_n15605));
  nor2 g15412(.a(new_n11596), .b(new_n1199), .O(new_n15606));
  inv1 g15413(.a(new_n15606), .O(new_n15607));
  nor2 g15414(.a(new_n15607), .b(new_n13306), .O(new_n15608));
  nor2 g15415(.a(new_n15608), .b(new_n15605), .O(new_n15609));
  inv1 g15416(.a(new_n15609), .O(new_n15610));
  nor2 g15417(.a(new_n15610), .b(new_n15603), .O(new_n15611));
  inv1 g15418(.a(new_n15603), .O(new_n15612));
  nor2 g15419(.a(new_n15609), .b(new_n15612), .O(new_n15613));
  nor2 g15420(.a(new_n15613), .b(new_n15611), .O(new_n15614));
  nor2 g15421(.a(new_n8026), .b(new_n1647), .O(new_n15615));
  inv1 g15422(.a(new_n15615), .O(new_n15616));
  nor2 g15423(.a(new_n4425), .b(new_n3870), .O(new_n15617));
  nor2 g15424(.a(new_n15617), .b(new_n15453), .O(new_n15618));
  inv1 g15425(.a(new_n15450), .O(new_n15619));
  nor2 g15426(.a(new_n4682), .b(new_n3870), .O(new_n15620));
  inv1 g15427(.a(new_n15620), .O(new_n15621));
  nor2 g15428(.a(new_n15621), .b(new_n15619), .O(new_n15622));
  nor2 g15429(.a(new_n15622), .b(new_n15618), .O(new_n15623));
  nor2 g15430(.a(new_n15623), .b(new_n15616), .O(new_n15624));
  inv1 g15431(.a(new_n15623), .O(new_n15625));
  nor2 g15432(.a(new_n15625), .b(new_n15615), .O(new_n15626));
  nor2 g15433(.a(new_n15626), .b(new_n15624), .O(new_n15627));
  nor2 g15434(.a(new_n15627), .b(new_n15614), .O(new_n15628));
  inv1 g15435(.a(new_n15614), .O(new_n15629));
  inv1 g15436(.a(new_n15627), .O(new_n15630));
  nor2 g15437(.a(new_n15630), .b(new_n15629), .O(new_n15631));
  nor2 g15438(.a(new_n15631), .b(new_n15628), .O(new_n15632));
  inv1 g15439(.a(new_n15632), .O(new_n15633));
  nor2 g15440(.a(new_n4366), .b(\a[37] ), .O(new_n15634));
  nor2 g15441(.a(new_n15634), .b(new_n15362), .O(new_n15635));
  inv1 g15442(.a(new_n15634), .O(new_n15636));
  nor2 g15443(.a(new_n15636), .b(new_n15361), .O(new_n15637));
  nor2 g15444(.a(new_n15637), .b(new_n15635), .O(new_n15638));
  nor2 g15445(.a(new_n15638), .b(new_n15633), .O(new_n15639));
  inv1 g15446(.a(new_n15638), .O(new_n15640));
  nor2 g15447(.a(new_n15640), .b(new_n15632), .O(new_n15641));
  nor2 g15448(.a(new_n15641), .b(new_n15639), .O(new_n15642));
  nor2 g15449(.a(new_n15642), .b(new_n15602), .O(new_n15643));
  inv1 g15450(.a(new_n15642), .O(new_n15644));
  nor2 g15451(.a(new_n15644), .b(new_n15601), .O(new_n15645));
  nor2 g15452(.a(new_n15645), .b(new_n15643), .O(new_n15646));
  inv1 g15453(.a(new_n15646), .O(new_n15647));
  nor2 g15454(.a(new_n6893), .b(new_n2184), .O(new_n15648));
  inv1 g15455(.a(new_n15648), .O(new_n15649));
  nor2 g15456(.a(new_n6274), .b(new_n2506), .O(new_n15650));
  nor2 g15457(.a(new_n15650), .b(new_n15384), .O(new_n15651));
  inv1 g15458(.a(new_n15381), .O(new_n15652));
  nor2 g15459(.a(new_n6570), .b(new_n2506), .O(new_n15653));
  inv1 g15460(.a(new_n15653), .O(new_n15654));
  nor2 g15461(.a(new_n15654), .b(new_n15652), .O(new_n15655));
  nor2 g15462(.a(new_n15655), .b(new_n15651), .O(new_n15656));
  nor2 g15463(.a(new_n15656), .b(new_n15649), .O(new_n15657));
  inv1 g15464(.a(new_n15656), .O(new_n15658));
  nor2 g15465(.a(new_n15658), .b(new_n15648), .O(new_n15659));
  nor2 g15466(.a(new_n15659), .b(new_n15657), .O(new_n15660));
  inv1 g15467(.a(new_n15660), .O(new_n15661));
  nor2 g15468(.a(new_n10895), .b(new_n699), .O(new_n15662));
  nor2 g15469(.a(new_n10468), .b(new_n800), .O(new_n15663));
  nor2 g15470(.a(new_n15663), .b(new_n15260), .O(new_n15664));
  inv1 g15471(.a(new_n15258), .O(new_n15665));
  nor2 g15472(.a(new_n10468), .b(new_n847), .O(new_n15666));
  inv1 g15473(.a(new_n15666), .O(new_n15667));
  nor2 g15474(.a(new_n15667), .b(new_n15665), .O(new_n15668));
  nor2 g15475(.a(new_n15668), .b(new_n15664), .O(new_n15669));
  inv1 g15476(.a(new_n15669), .O(new_n15670));
  nor2 g15477(.a(new_n15670), .b(new_n15662), .O(new_n15671));
  inv1 g15478(.a(new_n15662), .O(new_n15672));
  nor2 g15479(.a(new_n15669), .b(new_n15672), .O(new_n15673));
  nor2 g15480(.a(new_n15673), .b(new_n15671), .O(new_n15674));
  nor2 g15481(.a(new_n9873), .b(new_n941), .O(new_n15675));
  inv1 g15482(.a(new_n15675), .O(new_n15676));
  nor2 g15483(.a(new_n6958), .b(new_n2121), .O(new_n15677));
  nor2 g15484(.a(new_n9658), .b(new_n1086), .O(new_n15678));
  nor2 g15485(.a(new_n15678), .b(new_n15677), .O(new_n15679));
  nor2 g15486(.a(new_n9658), .b(new_n2121), .O(new_n15680));
  inv1 g15487(.a(new_n15680), .O(new_n15681));
  nor2 g15488(.a(new_n15681), .b(new_n13126), .O(new_n15682));
  nor2 g15489(.a(new_n15682), .b(new_n15679), .O(new_n15683));
  nor2 g15490(.a(new_n15683), .b(new_n15676), .O(new_n15684));
  inv1 g15491(.a(new_n15683), .O(new_n15685));
  nor2 g15492(.a(new_n15685), .b(new_n15675), .O(new_n15686));
  nor2 g15493(.a(new_n15686), .b(new_n15684), .O(new_n15687));
  nor2 g15494(.a(new_n15687), .b(new_n15674), .O(new_n15688));
  inv1 g15495(.a(new_n15674), .O(new_n15689));
  inv1 g15496(.a(new_n15687), .O(new_n15690));
  nor2 g15497(.a(new_n15690), .b(new_n15689), .O(new_n15691));
  nor2 g15498(.a(new_n15691), .b(new_n15688), .O(new_n15692));
  nor2 g15499(.a(new_n15692), .b(new_n15661), .O(new_n15693));
  inv1 g15500(.a(new_n15692), .O(new_n15694));
  nor2 g15501(.a(new_n15694), .b(new_n15660), .O(new_n15695));
  nor2 g15502(.a(new_n15695), .b(new_n15693), .O(new_n15696));
  inv1 g15503(.a(new_n15696), .O(new_n15697));
  nor2 g15504(.a(new_n15697), .b(new_n15647), .O(new_n15698));
  nor2 g15505(.a(new_n15696), .b(new_n15646), .O(new_n15699));
  nor2 g15506(.a(new_n15699), .b(new_n15698), .O(new_n15700));
  inv1 g15507(.a(new_n15700), .O(new_n15701));
  nor2 g15508(.a(new_n15701), .b(new_n15600), .O(new_n15702));
  nor2 g15509(.a(new_n15700), .b(new_n15599), .O(new_n15703));
  nor2 g15510(.a(new_n15703), .b(new_n15702), .O(new_n15704));
  nor2 g15511(.a(new_n15704), .b(new_n15568), .O(new_n15705));
  inv1 g15512(.a(new_n15568), .O(new_n15706));
  inv1 g15513(.a(new_n15704), .O(new_n15707));
  nor2 g15514(.a(new_n15707), .b(new_n15706), .O(new_n15708));
  nor2 g15515(.a(new_n15708), .b(new_n15705), .O(new_n15709));
  inv1 g15516(.a(new_n15709), .O(new_n15710));
  nor2 g15517(.a(new_n15479), .b(new_n15341), .O(new_n15711));
  inv1 g15518(.a(new_n15711), .O(new_n15712));
  nor2 g15519(.a(new_n15293), .b(new_n15287), .O(new_n15713));
  nor2 g15520(.a(new_n15282), .b(new_n15276), .O(new_n15714));
  nor2 g15521(.a(new_n15337), .b(new_n15334), .O(new_n15715));
  nor2 g15522(.a(new_n8476), .b(new_n1425), .O(new_n15716));
  inv1 g15523(.a(new_n15716), .O(new_n15717));
  nor2 g15524(.a(new_n8170), .b(new_n1493), .O(new_n15718));
  nor2 g15525(.a(new_n15718), .b(new_n15430), .O(new_n15719));
  nor2 g15526(.a(new_n8170), .b(new_n1736), .O(new_n15720));
  inv1 g15527(.a(new_n15720), .O(new_n15721));
  nor2 g15528(.a(new_n15721), .b(new_n14739), .O(new_n15722));
  nor2 g15529(.a(new_n15722), .b(new_n15719), .O(new_n15723));
  nor2 g15530(.a(new_n15723), .b(new_n15717), .O(new_n15724));
  inv1 g15531(.a(new_n15723), .O(new_n15725));
  nor2 g15532(.a(new_n15725), .b(new_n15716), .O(new_n15726));
  nor2 g15533(.a(new_n15726), .b(new_n15724), .O(new_n15727));
  nor2 g15534(.a(new_n5796), .b(new_n2826), .O(new_n15728));
  inv1 g15535(.a(new_n15728), .O(new_n15729));
  nor2 g15536(.a(new_n5178), .b(new_n3231), .O(new_n15730));
  nor2 g15537(.a(new_n15730), .b(new_n15397), .O(new_n15731));
  inv1 g15538(.a(new_n15395), .O(new_n15732));
  nor2 g15539(.a(new_n5393), .b(new_n3231), .O(new_n15733));
  inv1 g15540(.a(new_n15733), .O(new_n15734));
  nor2 g15541(.a(new_n15734), .b(new_n15732), .O(new_n15735));
  nor2 g15542(.a(new_n15735), .b(new_n15731), .O(new_n15736));
  nor2 g15543(.a(new_n15736), .b(new_n15729), .O(new_n15737));
  inv1 g15544(.a(new_n15736), .O(new_n15738));
  nor2 g15545(.a(new_n15738), .b(new_n15728), .O(new_n15739));
  nor2 g15546(.a(new_n15739), .b(new_n15737), .O(new_n15740));
  nor2 g15547(.a(new_n4954), .b(new_n3533), .O(new_n15741));
  inv1 g15548(.a(new_n15741), .O(new_n15742));
  nor2 g15549(.a(new_n8946), .b(new_n1297), .O(new_n15743));
  nor2 g15550(.a(new_n7294), .b(new_n1903), .O(new_n15744));
  nor2 g15551(.a(new_n15744), .b(new_n15743), .O(new_n15745));
  inv1 g15552(.a(new_n15743), .O(new_n15746));
  inv1 g15553(.a(new_n15744), .O(new_n15747));
  nor2 g15554(.a(new_n15747), .b(new_n15746), .O(new_n15748));
  nor2 g15555(.a(new_n15748), .b(new_n15745), .O(new_n15749));
  inv1 g15556(.a(new_n15749), .O(new_n15750));
  nor2 g15557(.a(new_n15750), .b(new_n15742), .O(new_n15751));
  nor2 g15558(.a(new_n15749), .b(new_n15741), .O(new_n15752));
  nor2 g15559(.a(new_n15752), .b(new_n15751), .O(new_n15753));
  inv1 g15560(.a(new_n15753), .O(new_n15754));
  nor2 g15561(.a(new_n15754), .b(new_n15740), .O(new_n15755));
  inv1 g15562(.a(new_n15740), .O(new_n15756));
  nor2 g15563(.a(new_n15753), .b(new_n15756), .O(new_n15757));
  nor2 g15564(.a(new_n15757), .b(new_n15755), .O(new_n15758));
  nor2 g15565(.a(new_n15758), .b(new_n15727), .O(new_n15759));
  inv1 g15566(.a(new_n15727), .O(new_n15760));
  inv1 g15567(.a(new_n15758), .O(new_n15761));
  nor2 g15568(.a(new_n15761), .b(new_n15760), .O(new_n15762));
  nor2 g15569(.a(new_n15762), .b(new_n15759), .O(new_n15763));
  nor2 g15570(.a(new_n15763), .b(new_n15715), .O(new_n15764));
  inv1 g15571(.a(new_n15715), .O(new_n15765));
  inv1 g15572(.a(new_n15763), .O(new_n15766));
  nor2 g15573(.a(new_n15766), .b(new_n15765), .O(new_n15767));
  nor2 g15574(.a(new_n15767), .b(new_n15764), .O(new_n15768));
  inv1 g15575(.a(new_n15768), .O(new_n15769));
  nor2 g15576(.a(new_n15769), .b(new_n15714), .O(new_n15770));
  inv1 g15577(.a(new_n15714), .O(new_n15771));
  nor2 g15578(.a(new_n15768), .b(new_n15771), .O(new_n15772));
  nor2 g15579(.a(new_n15772), .b(new_n15770), .O(new_n15773));
  inv1 g15580(.a(new_n15773), .O(new_n15774));
  nor2 g15581(.a(new_n15774), .b(new_n15713), .O(new_n15775));
  inv1 g15582(.a(new_n15713), .O(new_n15776));
  nor2 g15583(.a(new_n15773), .b(new_n15776), .O(new_n15777));
  nor2 g15584(.a(new_n15777), .b(new_n15775), .O(new_n15778));
  nor2 g15585(.a(new_n15778), .b(new_n15712), .O(new_n15779));
  inv1 g15586(.a(new_n15778), .O(new_n15780));
  nor2 g15587(.a(new_n15780), .b(new_n15711), .O(new_n15781));
  nor2 g15588(.a(new_n15781), .b(new_n15779), .O(new_n15782));
  inv1 g15589(.a(new_n15782), .O(new_n15783));
  nor2 g15590(.a(new_n15483), .b(new_n15297), .O(new_n15784));
  nor2 g15591(.a(new_n15784), .b(new_n15783), .O(new_n15785));
  inv1 g15592(.a(new_n15784), .O(new_n15786));
  nor2 g15593(.a(new_n15786), .b(new_n15782), .O(new_n15787));
  nor2 g15594(.a(new_n15787), .b(new_n15785), .O(new_n15788));
  inv1 g15595(.a(new_n15788), .O(new_n15789));
  nor2 g15596(.a(new_n15789), .b(new_n15710), .O(new_n15790));
  nor2 g15597(.a(new_n15788), .b(new_n15709), .O(new_n15791));
  nor2 g15598(.a(new_n15791), .b(new_n15790), .O(new_n15792));
  inv1 g15599(.a(new_n15792), .O(new_n15793));
  nor2 g15600(.a(new_n15793), .b(new_n15501), .O(new_n15794));
  inv1 g15601(.a(new_n15501), .O(new_n15795));
  nor2 g15602(.a(new_n15792), .b(new_n15795), .O(new_n15796));
  nor2 g15603(.a(new_n15796), .b(new_n15794), .O(new_n15797));
  inv1 g15604(.a(new_n15797), .O(new_n15798));
  nor2 g15605(.a(new_n15498), .b(new_n15490), .O(new_n15799));
  nor2 g15606(.a(new_n15799), .b(new_n15798), .O(new_n15800));
  inv1 g15607(.a(new_n15799), .O(new_n15801));
  nor2 g15608(.a(new_n15801), .b(new_n15797), .O(new_n15802));
  nor2 g15609(.a(new_n15802), .b(new_n15800), .O(new_n15803));
  inv1 g15610(.a(new_n15803), .O(\asquared[76] ));
  nor2 g15611(.a(new_n15790), .b(new_n15785), .O(new_n15805));
  nor2 g15612(.a(new_n15708), .b(new_n15567), .O(new_n15806));
  nor2 g15613(.a(new_n15702), .b(new_n15596), .O(new_n15807));
  nor2 g15614(.a(new_n15562), .b(new_n15519), .O(new_n15808));
  nor2 g15615(.a(new_n15557), .b(new_n15553), .O(new_n15809));
  nor2 g15616(.a(new_n15592), .b(new_n15589), .O(new_n15810));
  nor2 g15617(.a(new_n8476), .b(new_n1493), .O(new_n15811));
  nor2 g15618(.a(new_n15811), .b(new_n15441), .O(new_n15812));
  nor2 g15619(.a(new_n8946), .b(new_n1493), .O(new_n15813));
  inv1 g15620(.a(new_n15813), .O(new_n15814));
  nor2 g15621(.a(new_n15814), .b(new_n15717), .O(new_n15815));
  nor2 g15622(.a(new_n15815), .b(new_n15812), .O(new_n15816));
  nor2 g15623(.a(new_n15816), .b(new_n13005), .O(new_n15817));
  inv1 g15624(.a(new_n15816), .O(new_n15818));
  nor2 g15625(.a(new_n15818), .b(new_n13004), .O(new_n15819));
  nor2 g15626(.a(new_n15819), .b(new_n15817), .O(new_n15820));
  inv1 g15627(.a(new_n15820), .O(new_n15821));
  nor2 g15628(.a(new_n11596), .b(new_n613), .O(new_n15822));
  nor2 g15629(.a(new_n5971), .b(new_n2826), .O(new_n15823));
  nor2 g15630(.a(new_n5796), .b(new_n3057), .O(new_n15824));
  nor2 g15631(.a(new_n15824), .b(new_n15823), .O(new_n15825));
  nor2 g15632(.a(new_n5971), .b(new_n3057), .O(new_n15826));
  inv1 g15633(.a(new_n15826), .O(new_n15827));
  nor2 g15634(.a(new_n15827), .b(new_n15729), .O(new_n15828));
  nor2 g15635(.a(new_n15828), .b(new_n15825), .O(new_n15829));
  inv1 g15636(.a(new_n15829), .O(new_n15830));
  nor2 g15637(.a(new_n15830), .b(new_n15822), .O(new_n15831));
  inv1 g15638(.a(new_n15822), .O(new_n15832));
  nor2 g15639(.a(new_n15829), .b(new_n15832), .O(new_n15833));
  nor2 g15640(.a(new_n15833), .b(new_n15831), .O(new_n15834));
  nor2 g15641(.a(new_n9658), .b(new_n1199), .O(new_n15835));
  nor2 g15642(.a(new_n8170), .b(new_n1647), .O(new_n15836));
  nor2 g15643(.a(new_n15836), .b(new_n15835), .O(new_n15837));
  inv1 g15644(.a(new_n15835), .O(new_n15838));
  inv1 g15645(.a(new_n15836), .O(new_n15839));
  nor2 g15646(.a(new_n15839), .b(new_n15838), .O(new_n15840));
  nor2 g15647(.a(new_n15840), .b(new_n15837), .O(new_n15841));
  nor2 g15648(.a(new_n15841), .b(new_n15734), .O(new_n15842));
  inv1 g15649(.a(new_n15841), .O(new_n15843));
  nor2 g15650(.a(new_n15843), .b(new_n15733), .O(new_n15844));
  nor2 g15651(.a(new_n15844), .b(new_n15842), .O(new_n15845));
  nor2 g15652(.a(new_n15845), .b(new_n15834), .O(new_n15846));
  inv1 g15653(.a(new_n15834), .O(new_n15847));
  inv1 g15654(.a(new_n15845), .O(new_n15848));
  nor2 g15655(.a(new_n15848), .b(new_n15847), .O(new_n15849));
  nor2 g15656(.a(new_n15849), .b(new_n15846), .O(new_n15850));
  nor2 g15657(.a(new_n15850), .b(new_n15821), .O(new_n15851));
  inv1 g15658(.a(new_n15850), .O(new_n15852));
  nor2 g15659(.a(new_n15852), .b(new_n15820), .O(new_n15853));
  nor2 g15660(.a(new_n15853), .b(new_n15851), .O(new_n15854));
  inv1 g15661(.a(new_n15854), .O(new_n15855));
  nor2 g15662(.a(new_n15855), .b(new_n15810), .O(new_n15856));
  inv1 g15663(.a(new_n15810), .O(new_n15857));
  nor2 g15664(.a(new_n15854), .b(new_n15857), .O(new_n15858));
  nor2 g15665(.a(new_n15858), .b(new_n15856), .O(new_n15859));
  inv1 g15666(.a(new_n15859), .O(new_n15860));
  nor2 g15667(.a(new_n15860), .b(new_n15809), .O(new_n15861));
  inv1 g15668(.a(new_n15809), .O(new_n15862));
  nor2 g15669(.a(new_n15859), .b(new_n15862), .O(new_n15863));
  nor2 g15670(.a(new_n15863), .b(new_n15861), .O(new_n15864));
  inv1 g15671(.a(new_n15864), .O(new_n15865));
  nor2 g15672(.a(new_n15865), .b(new_n15808), .O(new_n15866));
  inv1 g15673(.a(new_n15808), .O(new_n15867));
  nor2 g15674(.a(new_n15864), .b(new_n15867), .O(new_n15868));
  nor2 g15675(.a(new_n15868), .b(new_n15866), .O(new_n15869));
  inv1 g15676(.a(new_n15869), .O(new_n15870));
  nor2 g15677(.a(new_n15870), .b(new_n15807), .O(new_n15871));
  inv1 g15678(.a(new_n15807), .O(new_n15872));
  nor2 g15679(.a(new_n15869), .b(new_n15872), .O(new_n15873));
  nor2 g15680(.a(new_n15873), .b(new_n15871), .O(new_n15874));
  inv1 g15681(.a(new_n15874), .O(new_n15875));
  nor2 g15682(.a(new_n15875), .b(new_n15806), .O(new_n15876));
  inv1 g15683(.a(new_n15806), .O(new_n15877));
  nor2 g15684(.a(new_n15874), .b(new_n15877), .O(new_n15878));
  nor2 g15685(.a(new_n15878), .b(new_n15876), .O(new_n15879));
  inv1 g15686(.a(new_n15879), .O(new_n15880));
  nor2 g15687(.a(new_n15781), .b(new_n15775), .O(new_n15881));
  inv1 g15688(.a(new_n15881), .O(new_n15882));
  nor2 g15689(.a(new_n15550), .b(new_n15544), .O(new_n15883));
  inv1 g15690(.a(new_n15883), .O(new_n15884));
  nor2 g15691(.a(new_n15581), .b(new_n15575), .O(new_n15885));
  inv1 g15692(.a(new_n15885), .O(new_n15886));
  nor2 g15693(.a(new_n15886), .b(new_n15884), .O(new_n15887));
  nor2 g15694(.a(new_n15885), .b(new_n15883), .O(new_n15888));
  nor2 g15695(.a(new_n15888), .b(new_n15887), .O(new_n15889));
  nor2 g15696(.a(new_n15536), .b(new_n15530), .O(new_n15890));
  inv1 g15697(.a(new_n15890), .O(new_n15891));
  nor2 g15698(.a(new_n15891), .b(new_n15889), .O(new_n15892));
  inv1 g15699(.a(new_n15889), .O(new_n15893));
  nor2 g15700(.a(new_n15890), .b(new_n15893), .O(new_n15894));
  nor2 g15701(.a(new_n15894), .b(new_n15892), .O(new_n15895));
  inv1 g15702(.a(new_n15895), .O(new_n15896));
  nor2 g15703(.a(new_n15698), .b(new_n15645), .O(new_n15897));
  nor2 g15704(.a(new_n15897), .b(new_n15896), .O(new_n15898));
  inv1 g15705(.a(new_n15897), .O(new_n15899));
  nor2 g15706(.a(new_n15899), .b(new_n15895), .O(new_n15900));
  nor2 g15707(.a(new_n15900), .b(new_n15898), .O(new_n15901));
  inv1 g15708(.a(new_n15901), .O(new_n15902));
  nor2 g15709(.a(new_n15751), .b(new_n15748), .O(new_n15903));
  inv1 g15710(.a(new_n15903), .O(new_n15904));
  nor2 g15711(.a(new_n15659), .b(new_n15651), .O(new_n15905));
  nor2 g15712(.a(new_n15905), .b(new_n15904), .O(new_n15906));
  inv1 g15713(.a(new_n15905), .O(new_n15907));
  nor2 g15714(.a(new_n15907), .b(new_n15903), .O(new_n15908));
  nor2 g15715(.a(new_n15908), .b(new_n15906), .O(new_n15909));
  nor2 g15716(.a(new_n15611), .b(new_n15605), .O(new_n15910));
  nor2 g15717(.a(new_n15910), .b(new_n15909), .O(new_n15911));
  inv1 g15718(.a(new_n15909), .O(new_n15912));
  inv1 g15719(.a(new_n15910), .O(new_n15913));
  nor2 g15720(.a(new_n15913), .b(new_n15912), .O(new_n15914));
  nor2 g15721(.a(new_n15914), .b(new_n15911), .O(new_n15915));
  inv1 g15722(.a(new_n15915), .O(new_n15916));
  nor2 g15723(.a(new_n11186), .b(new_n699), .O(new_n15917));
  nor2 g15724(.a(new_n15637), .b(new_n4366), .O(new_n15918));
  nor2 g15725(.a(new_n15918), .b(new_n15917), .O(new_n15919));
  inv1 g15726(.a(new_n15917), .O(new_n15920));
  inv1 g15727(.a(new_n15918), .O(new_n15921));
  nor2 g15728(.a(new_n15921), .b(new_n15920), .O(new_n15922));
  nor2 g15729(.a(new_n15922), .b(new_n15919), .O(new_n15923));
  inv1 g15730(.a(new_n15923), .O(new_n15924));
  nor2 g15731(.a(new_n15626), .b(new_n15618), .O(new_n15925));
  inv1 g15732(.a(new_n15925), .O(new_n15926));
  nor2 g15733(.a(new_n15926), .b(new_n15924), .O(new_n15927));
  nor2 g15734(.a(new_n15925), .b(new_n15923), .O(new_n15928));
  nor2 g15735(.a(new_n15928), .b(new_n15927), .O(new_n15929));
  inv1 g15736(.a(new_n15929), .O(new_n15930));
  nor2 g15737(.a(new_n15762), .b(new_n15757), .O(new_n15931));
  inv1 g15738(.a(new_n15931), .O(new_n15932));
  nor2 g15739(.a(new_n15932), .b(new_n15930), .O(new_n15933));
  nor2 g15740(.a(new_n15931), .b(new_n15929), .O(new_n15934));
  nor2 g15741(.a(new_n15934), .b(new_n15933), .O(new_n15935));
  inv1 g15742(.a(new_n15935), .O(new_n15936));
  nor2 g15743(.a(new_n15936), .b(new_n15916), .O(new_n15937));
  nor2 g15744(.a(new_n15935), .b(new_n15915), .O(new_n15938));
  nor2 g15745(.a(new_n15938), .b(new_n15937), .O(new_n15939));
  inv1 g15746(.a(new_n15939), .O(new_n15940));
  nor2 g15747(.a(new_n15940), .b(new_n15902), .O(new_n15941));
  nor2 g15748(.a(new_n15939), .b(new_n15901), .O(new_n15942));
  nor2 g15749(.a(new_n15942), .b(new_n15941), .O(new_n15943));
  nor2 g15750(.a(new_n15943), .b(new_n15882), .O(new_n15944));
  inv1 g15751(.a(new_n15943), .O(new_n15945));
  nor2 g15752(.a(new_n15945), .b(new_n15881), .O(new_n15946));
  nor2 g15753(.a(new_n15946), .b(new_n15944), .O(new_n15947));
  inv1 g15754(.a(new_n15947), .O(new_n15948));
  nor2 g15755(.a(new_n15770), .b(new_n15764), .O(new_n15949));
  inv1 g15756(.a(new_n15949), .O(new_n15950));
  nor2 g15757(.a(new_n15686), .b(new_n15679), .O(new_n15951));
  nor2 g15758(.a(new_n15671), .b(new_n15664), .O(new_n15952));
  nor2 g15759(.a(new_n15952), .b(new_n15951), .O(new_n15953));
  inv1 g15760(.a(new_n15951), .O(new_n15954));
  inv1 g15761(.a(new_n15952), .O(new_n15955));
  nor2 g15762(.a(new_n15955), .b(new_n15954), .O(new_n15956));
  nor2 g15763(.a(new_n15956), .b(new_n15953), .O(new_n15957));
  nor2 g15764(.a(new_n15739), .b(new_n15731), .O(new_n15958));
  nor2 g15765(.a(new_n15958), .b(new_n15957), .O(new_n15959));
  inv1 g15766(.a(new_n15957), .O(new_n15960));
  inv1 g15767(.a(new_n15958), .O(new_n15961));
  nor2 g15768(.a(new_n15961), .b(new_n15960), .O(new_n15962));
  nor2 g15769(.a(new_n15962), .b(new_n15959), .O(new_n15963));
  inv1 g15770(.a(new_n15963), .O(new_n15964));
  nor2 g15771(.a(new_n15695), .b(new_n15688), .O(new_n15965));
  inv1 g15772(.a(new_n15965), .O(new_n15966));
  nor2 g15773(.a(new_n15639), .b(new_n15628), .O(new_n15967));
  inv1 g15774(.a(new_n15967), .O(new_n15968));
  nor2 g15775(.a(new_n15968), .b(new_n15966), .O(new_n15969));
  nor2 g15776(.a(new_n15967), .b(new_n15965), .O(new_n15970));
  nor2 g15777(.a(new_n15970), .b(new_n15969), .O(new_n15971));
  inv1 g15778(.a(new_n15971), .O(new_n15972));
  nor2 g15779(.a(new_n15972), .b(new_n15964), .O(new_n15973));
  nor2 g15780(.a(new_n15971), .b(new_n15963), .O(new_n15974));
  nor2 g15781(.a(new_n15974), .b(new_n15973), .O(new_n15975));
  nor2 g15782(.a(new_n15975), .b(new_n15950), .O(new_n15976));
  inv1 g15783(.a(new_n15975), .O(new_n15977));
  nor2 g15784(.a(new_n15977), .b(new_n15949), .O(new_n15978));
  nor2 g15785(.a(new_n15978), .b(new_n15976), .O(new_n15979));
  inv1 g15786(.a(new_n15979), .O(new_n15980));
  nor2 g15787(.a(new_n15515), .b(new_n15509), .O(new_n15981));
  inv1 g15788(.a(new_n15981), .O(new_n15982));
  nor2 g15789(.a(new_n4425), .b(new_n4093), .O(new_n15983));
  inv1 g15790(.a(new_n15983), .O(new_n15984));
  nor2 g15791(.a(new_n7537), .b(new_n1903), .O(new_n15985));
  nor2 g15792(.a(new_n8026), .b(new_n1736), .O(new_n15986));
  nor2 g15793(.a(new_n15986), .b(new_n15985), .O(new_n15987));
  nor2 g15794(.a(new_n8026), .b(new_n1903), .O(new_n15988));
  inv1 g15795(.a(new_n15988), .O(new_n15989));
  nor2 g15796(.a(new_n15989), .b(new_n15431), .O(new_n15990));
  nor2 g15797(.a(new_n15990), .b(new_n15987), .O(new_n15991));
  nor2 g15798(.a(new_n15991), .b(new_n15984), .O(new_n15992));
  inv1 g15799(.a(new_n15991), .O(new_n15993));
  nor2 g15800(.a(new_n15993), .b(new_n15983), .O(new_n15994));
  nor2 g15801(.a(new_n15994), .b(new_n15992), .O(new_n15995));
  inv1 g15802(.a(new_n15995), .O(new_n15996));
  nor2 g15803(.a(new_n6893), .b(new_n2433), .O(new_n15997));
  nor2 g15804(.a(new_n6274), .b(new_n2660), .O(new_n15998));
  nor2 g15805(.a(new_n15998), .b(new_n15653), .O(new_n15999));
  inv1 g15806(.a(new_n15650), .O(new_n16000));
  nor2 g15807(.a(new_n6570), .b(new_n2660), .O(new_n16001));
  inv1 g15808(.a(new_n16001), .O(new_n16002));
  nor2 g15809(.a(new_n16002), .b(new_n16000), .O(new_n16003));
  nor2 g15810(.a(new_n16003), .b(new_n15999), .O(new_n16004));
  inv1 g15811(.a(new_n16004), .O(new_n16005));
  nor2 g15812(.a(new_n16005), .b(new_n15997), .O(new_n16006));
  inv1 g15813(.a(new_n15997), .O(new_n16007));
  nor2 g15814(.a(new_n16004), .b(new_n16007), .O(new_n16008));
  nor2 g15815(.a(new_n16008), .b(new_n16006), .O(new_n16009));
  nor2 g15816(.a(new_n5178), .b(new_n3533), .O(new_n16010));
  inv1 g15817(.a(new_n16010), .O(new_n16011));
  nor2 g15818(.a(new_n4954), .b(new_n3722), .O(new_n16012));
  nor2 g15819(.a(new_n16012), .b(new_n15620), .O(new_n16013));
  nor2 g15820(.a(new_n4954), .b(new_n3870), .O(new_n16014));
  inv1 g15821(.a(new_n16014), .O(new_n16015));
  nor2 g15822(.a(new_n16015), .b(new_n15454), .O(new_n16016));
  nor2 g15823(.a(new_n16016), .b(new_n16013), .O(new_n16017));
  nor2 g15824(.a(new_n16017), .b(new_n16011), .O(new_n16018));
  inv1 g15825(.a(new_n16017), .O(new_n16019));
  nor2 g15826(.a(new_n16019), .b(new_n16010), .O(new_n16020));
  nor2 g15827(.a(new_n16020), .b(new_n16018), .O(new_n16021));
  nor2 g15828(.a(new_n16021), .b(new_n16009), .O(new_n16022));
  inv1 g15829(.a(new_n16009), .O(new_n16023));
  inv1 g15830(.a(new_n16021), .O(new_n16024));
  nor2 g15831(.a(new_n16024), .b(new_n16023), .O(new_n16025));
  nor2 g15832(.a(new_n16025), .b(new_n16022), .O(new_n16026));
  nor2 g15833(.a(new_n16026), .b(new_n15996), .O(new_n16027));
  inv1 g15834(.a(new_n16026), .O(new_n16028));
  nor2 g15835(.a(new_n16028), .b(new_n15995), .O(new_n16029));
  nor2 g15836(.a(new_n16029), .b(new_n16027), .O(new_n16030));
  nor2 g15837(.a(new_n16030), .b(new_n15982), .O(new_n16031));
  inv1 g15838(.a(new_n16030), .O(new_n16032));
  nor2 g15839(.a(new_n16032), .b(new_n15981), .O(new_n16033));
  nor2 g15840(.a(new_n16033), .b(new_n16031), .O(new_n16034));
  inv1 g15841(.a(new_n16034), .O(new_n16035));
  nor2 g15842(.a(new_n9873), .b(new_n1086), .O(new_n16036));
  inv1 g15843(.a(new_n16036), .O(new_n16037));
  nor2 g15844(.a(new_n7294), .b(new_n2121), .O(new_n16038));
  nor2 g15845(.a(new_n6958), .b(new_n2184), .O(new_n16039));
  nor2 g15846(.a(new_n16039), .b(new_n16038), .O(new_n16040));
  inv1 g15847(.a(new_n15677), .O(new_n16041));
  nor2 g15848(.a(new_n7294), .b(new_n2184), .O(new_n16042));
  inv1 g15849(.a(new_n16042), .O(new_n16043));
  nor2 g15850(.a(new_n16043), .b(new_n16041), .O(new_n16044));
  nor2 g15851(.a(new_n16044), .b(new_n16040), .O(new_n16045));
  nor2 g15852(.a(new_n16045), .b(new_n16037), .O(new_n16046));
  inv1 g15853(.a(new_n16045), .O(new_n16047));
  nor2 g15854(.a(new_n16047), .b(new_n16036), .O(new_n16048));
  nor2 g15855(.a(new_n16048), .b(new_n16046), .O(new_n16049));
  nor2 g15856(.a(new_n10895), .b(new_n800), .O(new_n16050));
  inv1 g15857(.a(new_n16050), .O(new_n16051));
  nor2 g15858(.a(new_n10320), .b(new_n941), .O(new_n16052));
  nor2 g15859(.a(new_n16052), .b(new_n15666), .O(new_n16053));
  nor2 g15860(.a(new_n10468), .b(new_n941), .O(new_n16054));
  inv1 g15861(.a(new_n16054), .O(new_n16055));
  nor2 g15862(.a(new_n16055), .b(new_n15261), .O(new_n16056));
  nor2 g15863(.a(new_n16056), .b(new_n16053), .O(new_n16057));
  nor2 g15864(.a(new_n16057), .b(new_n16051), .O(new_n16058));
  inv1 g15865(.a(new_n16057), .O(new_n16059));
  nor2 g15866(.a(new_n16059), .b(new_n16050), .O(new_n16060));
  nor2 g15867(.a(new_n16060), .b(new_n16058), .O(new_n16061));
  nor2 g15868(.a(new_n15726), .b(new_n15719), .O(new_n16062));
  inv1 g15869(.a(new_n16062), .O(new_n16063));
  nor2 g15870(.a(new_n16063), .b(new_n16061), .O(new_n16064));
  inv1 g15871(.a(new_n16061), .O(new_n16065));
  nor2 g15872(.a(new_n16062), .b(new_n16065), .O(new_n16066));
  nor2 g15873(.a(new_n16066), .b(new_n16064), .O(new_n16067));
  inv1 g15874(.a(new_n16067), .O(new_n16068));
  nor2 g15875(.a(new_n16068), .b(new_n16049), .O(new_n16069));
  inv1 g15876(.a(new_n16049), .O(new_n16070));
  nor2 g15877(.a(new_n16067), .b(new_n16070), .O(new_n16071));
  nor2 g15878(.a(new_n16071), .b(new_n16069), .O(new_n16072));
  inv1 g15879(.a(new_n16072), .O(new_n16073));
  nor2 g15880(.a(new_n16073), .b(new_n16035), .O(new_n16074));
  nor2 g15881(.a(new_n16072), .b(new_n16034), .O(new_n16075));
  nor2 g15882(.a(new_n16075), .b(new_n16074), .O(new_n16076));
  inv1 g15883(.a(new_n16076), .O(new_n16077));
  nor2 g15884(.a(new_n16077), .b(new_n15980), .O(new_n16078));
  nor2 g15885(.a(new_n16076), .b(new_n15979), .O(new_n16079));
  nor2 g15886(.a(new_n16079), .b(new_n16078), .O(new_n16080));
  inv1 g15887(.a(new_n16080), .O(new_n16081));
  nor2 g15888(.a(new_n16081), .b(new_n15948), .O(new_n16082));
  nor2 g15889(.a(new_n16080), .b(new_n15947), .O(new_n16083));
  nor2 g15890(.a(new_n16083), .b(new_n16082), .O(new_n16084));
  inv1 g15891(.a(new_n16084), .O(new_n16085));
  nor2 g15892(.a(new_n16085), .b(new_n15880), .O(new_n16086));
  nor2 g15893(.a(new_n16084), .b(new_n15879), .O(new_n16087));
  nor2 g15894(.a(new_n16087), .b(new_n16086), .O(new_n16088));
  inv1 g15895(.a(new_n16088), .O(new_n16089));
  nor2 g15896(.a(new_n16089), .b(new_n15805), .O(new_n16090));
  inv1 g15897(.a(new_n15805), .O(new_n16091));
  nor2 g15898(.a(new_n16088), .b(new_n16091), .O(new_n16092));
  nor2 g15899(.a(new_n16092), .b(new_n16090), .O(new_n16093));
  inv1 g15900(.a(new_n16093), .O(new_n16094));
  nor2 g15901(.a(new_n15800), .b(new_n15796), .O(new_n16095));
  nor2 g15902(.a(new_n16095), .b(new_n16094), .O(new_n16096));
  inv1 g15903(.a(new_n16095), .O(new_n16097));
  nor2 g15904(.a(new_n16097), .b(new_n16093), .O(new_n16098));
  nor2 g15905(.a(new_n16098), .b(new_n16096), .O(new_n16099));
  inv1 g15906(.a(new_n16099), .O(\asquared[77] ));
  nor2 g15907(.a(new_n16086), .b(new_n15876), .O(new_n16101));
  nor2 g15908(.a(new_n16082), .b(new_n15946), .O(new_n16102));
  nor2 g15909(.a(new_n16078), .b(new_n15978), .O(new_n16103));
  nor2 g15910(.a(new_n15941), .b(new_n15898), .O(new_n16104));
  nor2 g15911(.a(new_n15937), .b(new_n15933), .O(new_n16105));
  nor2 g15912(.a(new_n15973), .b(new_n15970), .O(new_n16106));
  nor2 g15913(.a(new_n10895), .b(new_n847), .O(new_n16107));
  inv1 g15914(.a(new_n16107), .O(new_n16108));
  nor2 g15915(.a(new_n5796), .b(new_n3231), .O(new_n16109));
  nor2 g15916(.a(new_n16109), .b(new_n15826), .O(new_n16110));
  inv1 g15917(.a(new_n15824), .O(new_n16111));
  nor2 g15918(.a(new_n5971), .b(new_n3231), .O(new_n16112));
  inv1 g15919(.a(new_n16112), .O(new_n16113));
  nor2 g15920(.a(new_n16113), .b(new_n16111), .O(new_n16114));
  nor2 g15921(.a(new_n16114), .b(new_n16110), .O(new_n16115));
  nor2 g15922(.a(new_n16115), .b(new_n16108), .O(new_n16116));
  inv1 g15923(.a(new_n16115), .O(new_n16117));
  nor2 g15924(.a(new_n16117), .b(new_n16107), .O(new_n16118));
  nor2 g15925(.a(new_n16118), .b(new_n16116), .O(new_n16119));
  nor2 g15926(.a(new_n8476), .b(new_n1647), .O(new_n16120));
  nor2 g15927(.a(new_n16120), .b(new_n15720), .O(new_n16121));
  nor2 g15928(.a(new_n15839), .b(new_n15031), .O(new_n16122));
  nor2 g15929(.a(new_n16122), .b(new_n16121), .O(new_n16123));
  nor2 g15930(.a(new_n16123), .b(new_n15989), .O(new_n16124));
  inv1 g15931(.a(new_n16123), .O(new_n16125));
  nor2 g15932(.a(new_n16125), .b(new_n15988), .O(new_n16126));
  nor2 g15933(.a(new_n16126), .b(new_n16124), .O(new_n16127));
  nor2 g15934(.a(new_n5393), .b(new_n3533), .O(new_n16128));
  inv1 g15935(.a(new_n16128), .O(new_n16129));
  nor2 g15936(.a(new_n7537), .b(new_n2121), .O(new_n16130));
  nor2 g15937(.a(new_n16130), .b(new_n15813), .O(new_n16131));
  inv1 g15938(.a(new_n16130), .O(new_n16132));
  nor2 g15939(.a(new_n16132), .b(new_n15814), .O(new_n16133));
  nor2 g15940(.a(new_n16133), .b(new_n16131), .O(new_n16134));
  inv1 g15941(.a(new_n16134), .O(new_n16135));
  nor2 g15942(.a(new_n16135), .b(new_n16129), .O(new_n16136));
  nor2 g15943(.a(new_n16134), .b(new_n16128), .O(new_n16137));
  nor2 g15944(.a(new_n16137), .b(new_n16136), .O(new_n16138));
  inv1 g15945(.a(new_n16138), .O(new_n16139));
  nor2 g15946(.a(new_n16139), .b(new_n16127), .O(new_n16140));
  inv1 g15947(.a(new_n16127), .O(new_n16141));
  nor2 g15948(.a(new_n16138), .b(new_n16141), .O(new_n16142));
  nor2 g15949(.a(new_n16142), .b(new_n16140), .O(new_n16143));
  nor2 g15950(.a(new_n16143), .b(new_n16119), .O(new_n16144));
  inv1 g15951(.a(new_n16119), .O(new_n16145));
  inv1 g15952(.a(new_n16143), .O(new_n16146));
  nor2 g15953(.a(new_n16146), .b(new_n16145), .O(new_n16147));
  nor2 g15954(.a(new_n16147), .b(new_n16144), .O(new_n16148));
  nor2 g15955(.a(new_n16148), .b(new_n16106), .O(new_n16149));
  inv1 g15956(.a(new_n16106), .O(new_n16150));
  inv1 g15957(.a(new_n16148), .O(new_n16151));
  nor2 g15958(.a(new_n16151), .b(new_n16150), .O(new_n16152));
  nor2 g15959(.a(new_n16152), .b(new_n16149), .O(new_n16153));
  inv1 g15960(.a(new_n16153), .O(new_n16154));
  nor2 g15961(.a(new_n16154), .b(new_n16105), .O(new_n16155));
  inv1 g15962(.a(new_n16105), .O(new_n16156));
  nor2 g15963(.a(new_n16153), .b(new_n16156), .O(new_n16157));
  nor2 g15964(.a(new_n16157), .b(new_n16155), .O(new_n16158));
  inv1 g15965(.a(new_n16158), .O(new_n16159));
  nor2 g15966(.a(new_n16159), .b(new_n16104), .O(new_n16160));
  inv1 g15967(.a(new_n16104), .O(new_n16161));
  nor2 g15968(.a(new_n16158), .b(new_n16161), .O(new_n16162));
  nor2 g15969(.a(new_n16162), .b(new_n16160), .O(new_n16163));
  inv1 g15970(.a(new_n16163), .O(new_n16164));
  nor2 g15971(.a(new_n16164), .b(new_n16103), .O(new_n16165));
  inv1 g15972(.a(new_n16103), .O(new_n16166));
  nor2 g15973(.a(new_n16163), .b(new_n16166), .O(new_n16167));
  nor2 g15974(.a(new_n16167), .b(new_n16165), .O(new_n16168));
  inv1 g15975(.a(new_n16168), .O(new_n16169));
  nor2 g15976(.a(new_n16169), .b(new_n16102), .O(new_n16170));
  inv1 g15977(.a(new_n16102), .O(new_n16171));
  nor2 g15978(.a(new_n16168), .b(new_n16171), .O(new_n16172));
  nor2 g15979(.a(new_n16172), .b(new_n16170), .O(new_n16173));
  inv1 g15980(.a(new_n16173), .O(new_n16174));
  nor2 g15981(.a(new_n15871), .b(new_n15866), .O(new_n16175));
  inv1 g15982(.a(new_n16175), .O(new_n16176));
  nor2 g15983(.a(new_n15962), .b(new_n15956), .O(new_n16177));
  inv1 g15984(.a(new_n16177), .O(new_n16178));
  nor2 g15985(.a(new_n10320), .b(new_n1086), .O(new_n16179));
  nor2 g15986(.a(new_n16179), .b(new_n16054), .O(new_n16180));
  inv1 g15987(.a(new_n16052), .O(new_n16181));
  nor2 g15988(.a(new_n10468), .b(new_n1086), .O(new_n16182));
  inv1 g15989(.a(new_n16182), .O(new_n16183));
  nor2 g15990(.a(new_n16183), .b(new_n16181), .O(new_n16184));
  nor2 g15991(.a(new_n16184), .b(new_n16180), .O(new_n16185));
  inv1 g15992(.a(new_n16185), .O(new_n16186));
  nor2 g15993(.a(new_n15994), .b(new_n15987), .O(new_n16187));
  inv1 g15994(.a(new_n16187), .O(new_n16188));
  nor2 g15995(.a(new_n16188), .b(new_n16186), .O(new_n16189));
  nor2 g15996(.a(new_n16187), .b(new_n16185), .O(new_n16190));
  nor2 g15997(.a(new_n16190), .b(new_n16189), .O(new_n16191));
  nor2 g15998(.a(new_n16191), .b(new_n16178), .O(new_n16192));
  inv1 g15999(.a(new_n16191), .O(new_n16193));
  nor2 g16000(.a(new_n16193), .b(new_n16177), .O(new_n16194));
  nor2 g16001(.a(new_n16194), .b(new_n16192), .O(new_n16195));
  nor2 g16002(.a(new_n15914), .b(new_n15908), .O(new_n16196));
  inv1 g16003(.a(new_n16196), .O(new_n16197));
  nor2 g16004(.a(new_n16197), .b(new_n16195), .O(new_n16198));
  inv1 g16005(.a(new_n16195), .O(new_n16199));
  nor2 g16006(.a(new_n16196), .b(new_n16199), .O(new_n16200));
  nor2 g16007(.a(new_n16200), .b(new_n16198), .O(new_n16201));
  inv1 g16008(.a(new_n16201), .O(new_n16202));
  nor2 g16009(.a(new_n16074), .b(new_n16033), .O(new_n16203));
  nor2 g16010(.a(new_n16203), .b(new_n16202), .O(new_n16204));
  inv1 g16011(.a(new_n16203), .O(new_n16205));
  nor2 g16012(.a(new_n16205), .b(new_n16201), .O(new_n16206));
  nor2 g16013(.a(new_n16206), .b(new_n16204), .O(new_n16207));
  inv1 g16014(.a(new_n16207), .O(new_n16208));
  nor2 g16015(.a(new_n15819), .b(new_n15812), .O(new_n16209));
  nor2 g16016(.a(new_n16006), .b(new_n15999), .O(new_n16210));
  nor2 g16017(.a(new_n16210), .b(new_n16209), .O(new_n16211));
  inv1 g16018(.a(new_n16209), .O(new_n16212));
  inv1 g16019(.a(new_n16210), .O(new_n16213));
  nor2 g16020(.a(new_n16213), .b(new_n16212), .O(new_n16214));
  nor2 g16021(.a(new_n16214), .b(new_n16211), .O(new_n16215));
  nor2 g16022(.a(new_n15831), .b(new_n15825), .O(new_n16216));
  nor2 g16023(.a(new_n16216), .b(new_n16215), .O(new_n16217));
  inv1 g16024(.a(new_n16215), .O(new_n16218));
  inv1 g16025(.a(new_n16216), .O(new_n16219));
  nor2 g16026(.a(new_n16219), .b(new_n16218), .O(new_n16220));
  nor2 g16027(.a(new_n16220), .b(new_n16217), .O(new_n16221));
  inv1 g16028(.a(new_n16221), .O(new_n16222));
  nor2 g16029(.a(new_n16060), .b(new_n16053), .O(new_n16223));
  nor2 g16030(.a(new_n16048), .b(new_n16040), .O(new_n16224));
  nor2 g16031(.a(new_n16224), .b(new_n16223), .O(new_n16225));
  inv1 g16032(.a(new_n16223), .O(new_n16226));
  inv1 g16033(.a(new_n16224), .O(new_n16227));
  nor2 g16034(.a(new_n16227), .b(new_n16226), .O(new_n16228));
  nor2 g16035(.a(new_n16228), .b(new_n16225), .O(new_n16229));
  nor2 g16036(.a(new_n15844), .b(new_n15837), .O(new_n16230));
  nor2 g16037(.a(new_n16230), .b(new_n16229), .O(new_n16231));
  inv1 g16038(.a(new_n16229), .O(new_n16232));
  inv1 g16039(.a(new_n16230), .O(new_n16233));
  nor2 g16040(.a(new_n16233), .b(new_n16232), .O(new_n16234));
  nor2 g16041(.a(new_n16234), .b(new_n16231), .O(new_n16235));
  nor2 g16042(.a(new_n15853), .b(new_n15846), .O(new_n16236));
  inv1 g16043(.a(new_n16236), .O(new_n16237));
  nor2 g16044(.a(new_n16237), .b(new_n16235), .O(new_n16238));
  inv1 g16045(.a(new_n16235), .O(new_n16239));
  nor2 g16046(.a(new_n16236), .b(new_n16239), .O(new_n16240));
  nor2 g16047(.a(new_n16240), .b(new_n16238), .O(new_n16241));
  inv1 g16048(.a(new_n16241), .O(new_n16242));
  nor2 g16049(.a(new_n16242), .b(new_n16222), .O(new_n16243));
  nor2 g16050(.a(new_n16241), .b(new_n16221), .O(new_n16244));
  nor2 g16051(.a(new_n16244), .b(new_n16243), .O(new_n16245));
  inv1 g16052(.a(new_n16245), .O(new_n16246));
  nor2 g16053(.a(new_n16246), .b(new_n16208), .O(new_n16247));
  nor2 g16054(.a(new_n16245), .b(new_n16207), .O(new_n16248));
  nor2 g16055(.a(new_n16248), .b(new_n16247), .O(new_n16249));
  nor2 g16056(.a(new_n16249), .b(new_n16176), .O(new_n16250));
  inv1 g16057(.a(new_n16249), .O(new_n16251));
  nor2 g16058(.a(new_n16251), .b(new_n16175), .O(new_n16252));
  nor2 g16059(.a(new_n16252), .b(new_n16250), .O(new_n16253));
  inv1 g16060(.a(new_n16253), .O(new_n16254));
  nor2 g16061(.a(new_n15927), .b(new_n15922), .O(new_n16255));
  inv1 g16062(.a(new_n16255), .O(new_n16256));
  nor2 g16063(.a(new_n16069), .b(new_n16064), .O(new_n16257));
  inv1 g16064(.a(new_n16257), .O(new_n16258));
  nor2 g16065(.a(new_n16258), .b(new_n16256), .O(new_n16259));
  nor2 g16066(.a(new_n16257), .b(new_n16255), .O(new_n16260));
  nor2 g16067(.a(new_n16260), .b(new_n16259), .O(new_n16261));
  nor2 g16068(.a(new_n16029), .b(new_n16022), .O(new_n16262));
  inv1 g16069(.a(new_n16262), .O(new_n16263));
  nor2 g16070(.a(new_n16263), .b(new_n16261), .O(new_n16264));
  inv1 g16071(.a(new_n16261), .O(new_n16265));
  nor2 g16072(.a(new_n16262), .b(new_n16265), .O(new_n16266));
  nor2 g16073(.a(new_n16266), .b(new_n16264), .O(new_n16267));
  nor2 g16074(.a(new_n15861), .b(new_n15856), .O(new_n16268));
  inv1 g16075(.a(new_n16268), .O(new_n16269));
  nor2 g16076(.a(new_n16269), .b(new_n16267), .O(new_n16270));
  inv1 g16077(.a(new_n16267), .O(new_n16271));
  nor2 g16078(.a(new_n16268), .b(new_n16271), .O(new_n16272));
  nor2 g16079(.a(new_n16272), .b(new_n16270), .O(new_n16273));
  inv1 g16080(.a(new_n16273), .O(new_n16274));
  nor2 g16081(.a(new_n15894), .b(new_n15888), .O(new_n16275));
  inv1 g16082(.a(new_n16275), .O(new_n16276));
  nor2 g16083(.a(new_n5178), .b(new_n3722), .O(new_n16277));
  inv1 g16084(.a(new_n16277), .O(new_n16278));
  nor2 g16085(.a(new_n4682), .b(new_n4093), .O(new_n16279));
  nor2 g16086(.a(new_n16279), .b(new_n16014), .O(new_n16280));
  nor2 g16087(.a(new_n4954), .b(new_n4093), .O(new_n16281));
  inv1 g16088(.a(new_n16281), .O(new_n16282));
  nor2 g16089(.a(new_n16282), .b(new_n15621), .O(new_n16283));
  nor2 g16090(.a(new_n16283), .b(new_n16280), .O(new_n16284));
  nor2 g16091(.a(new_n16284), .b(new_n16278), .O(new_n16285));
  inv1 g16092(.a(new_n16284), .O(new_n16286));
  nor2 g16093(.a(new_n16286), .b(new_n16277), .O(new_n16287));
  nor2 g16094(.a(new_n16287), .b(new_n16285), .O(new_n16288));
  nor2 g16095(.a(new_n11596), .b(new_n699), .O(new_n16289));
  nor2 g16096(.a(new_n6274), .b(new_n2826), .O(new_n16290));
  nor2 g16097(.a(new_n16290), .b(new_n16289), .O(new_n16291));
  nor2 g16098(.a(new_n11596), .b(new_n2826), .O(new_n16292));
  inv1 g16099(.a(new_n16292), .O(new_n16293));
  nor2 g16100(.a(new_n16293), .b(new_n9110), .O(new_n16294));
  nor2 g16101(.a(new_n16294), .b(new_n16291), .O(new_n16295));
  nor2 g16102(.a(new_n16295), .b(new_n16002), .O(new_n16296));
  inv1 g16103(.a(new_n16295), .O(new_n16297));
  nor2 g16104(.a(new_n16297), .b(new_n16001), .O(new_n16298));
  nor2 g16105(.a(new_n16298), .b(new_n16296), .O(new_n16299));
  nor2 g16106(.a(new_n16299), .b(new_n16288), .O(new_n16300));
  inv1 g16107(.a(new_n16288), .O(new_n16301));
  inv1 g16108(.a(new_n16299), .O(new_n16302));
  nor2 g16109(.a(new_n16302), .b(new_n16301), .O(new_n16303));
  nor2 g16110(.a(new_n16303), .b(new_n16300), .O(new_n16304));
  inv1 g16111(.a(new_n16304), .O(new_n16305));
  nor2 g16112(.a(new_n11186), .b(new_n800), .O(new_n16306));
  inv1 g16113(.a(new_n16306), .O(new_n16307));
  nor2 g16114(.a(new_n4425), .b(\a[38] ), .O(new_n16308));
  nor2 g16115(.a(new_n16308), .b(new_n16307), .O(new_n16309));
  inv1 g16116(.a(new_n16308), .O(new_n16310));
  nor2 g16117(.a(new_n16310), .b(new_n16306), .O(new_n16311));
  nor2 g16118(.a(new_n16311), .b(new_n16309), .O(new_n16312));
  nor2 g16119(.a(new_n16312), .b(new_n16305), .O(new_n16313));
  inv1 g16120(.a(new_n16312), .O(new_n16314));
  nor2 g16121(.a(new_n16314), .b(new_n16304), .O(new_n16315));
  nor2 g16122(.a(new_n16315), .b(new_n16313), .O(new_n16316));
  nor2 g16123(.a(new_n16316), .b(new_n16276), .O(new_n16317));
  inv1 g16124(.a(new_n16316), .O(new_n16318));
  nor2 g16125(.a(new_n16318), .b(new_n16275), .O(new_n16319));
  nor2 g16126(.a(new_n16319), .b(new_n16317), .O(new_n16320));
  inv1 g16127(.a(new_n16320), .O(new_n16321));
  nor2 g16128(.a(new_n6958), .b(new_n2433), .O(new_n16322));
  nor2 g16129(.a(new_n6893), .b(new_n2506), .O(new_n16323));
  nor2 g16130(.a(new_n16323), .b(new_n16322), .O(new_n16324));
  nor2 g16131(.a(new_n6958), .b(new_n2506), .O(new_n16325));
  inv1 g16132(.a(new_n16325), .O(new_n16326));
  nor2 g16133(.a(new_n16326), .b(new_n16007), .O(new_n16327));
  nor2 g16134(.a(new_n16327), .b(new_n16324), .O(new_n16328));
  nor2 g16135(.a(new_n16328), .b(new_n16043), .O(new_n16329));
  inv1 g16136(.a(new_n16328), .O(new_n16330));
  nor2 g16137(.a(new_n16330), .b(new_n16042), .O(new_n16331));
  nor2 g16138(.a(new_n16331), .b(new_n16329), .O(new_n16332));
  nor2 g16139(.a(new_n9873), .b(new_n1199), .O(new_n16333));
  inv1 g16140(.a(new_n16333), .O(new_n16334));
  nor2 g16141(.a(new_n9658), .b(new_n1297), .O(new_n16335));
  nor2 g16142(.a(new_n9156), .b(new_n1425), .O(new_n16336));
  nor2 g16143(.a(new_n16336), .b(new_n16335), .O(new_n16337));
  nor2 g16144(.a(new_n9658), .b(new_n1425), .O(new_n16338));
  inv1 g16145(.a(new_n16338), .O(new_n16339));
  nor2 g16146(.a(new_n16339), .b(new_n13005), .O(new_n16340));
  nor2 g16147(.a(new_n16340), .b(new_n16337), .O(new_n16341));
  nor2 g16148(.a(new_n16341), .b(new_n16334), .O(new_n16342));
  inv1 g16149(.a(new_n16341), .O(new_n16343));
  nor2 g16150(.a(new_n16343), .b(new_n16333), .O(new_n16344));
  nor2 g16151(.a(new_n16344), .b(new_n16342), .O(new_n16345));
  nor2 g16152(.a(new_n16020), .b(new_n16013), .O(new_n16346));
  inv1 g16153(.a(new_n16346), .O(new_n16347));
  nor2 g16154(.a(new_n16347), .b(new_n16345), .O(new_n16348));
  inv1 g16155(.a(new_n16345), .O(new_n16349));
  nor2 g16156(.a(new_n16346), .b(new_n16349), .O(new_n16350));
  nor2 g16157(.a(new_n16350), .b(new_n16348), .O(new_n16351));
  inv1 g16158(.a(new_n16351), .O(new_n16352));
  nor2 g16159(.a(new_n16352), .b(new_n16332), .O(new_n16353));
  inv1 g16160(.a(new_n16332), .O(new_n16354));
  nor2 g16161(.a(new_n16351), .b(new_n16354), .O(new_n16355));
  nor2 g16162(.a(new_n16355), .b(new_n16353), .O(new_n16356));
  inv1 g16163(.a(new_n16356), .O(new_n16357));
  nor2 g16164(.a(new_n16357), .b(new_n16321), .O(new_n16358));
  nor2 g16165(.a(new_n16356), .b(new_n16320), .O(new_n16359));
  nor2 g16166(.a(new_n16359), .b(new_n16358), .O(new_n16360));
  inv1 g16167(.a(new_n16360), .O(new_n16361));
  nor2 g16168(.a(new_n16361), .b(new_n16274), .O(new_n16362));
  nor2 g16169(.a(new_n16360), .b(new_n16273), .O(new_n16363));
  nor2 g16170(.a(new_n16363), .b(new_n16362), .O(new_n16364));
  inv1 g16171(.a(new_n16364), .O(new_n16365));
  nor2 g16172(.a(new_n16365), .b(new_n16254), .O(new_n16366));
  nor2 g16173(.a(new_n16364), .b(new_n16253), .O(new_n16367));
  nor2 g16174(.a(new_n16367), .b(new_n16366), .O(new_n16368));
  inv1 g16175(.a(new_n16368), .O(new_n16369));
  nor2 g16176(.a(new_n16369), .b(new_n16174), .O(new_n16370));
  nor2 g16177(.a(new_n16368), .b(new_n16173), .O(new_n16371));
  nor2 g16178(.a(new_n16371), .b(new_n16370), .O(new_n16372));
  inv1 g16179(.a(new_n16372), .O(new_n16373));
  nor2 g16180(.a(new_n16373), .b(new_n16101), .O(new_n16374));
  inv1 g16181(.a(new_n16101), .O(new_n16375));
  nor2 g16182(.a(new_n16372), .b(new_n16375), .O(new_n16376));
  nor2 g16183(.a(new_n16376), .b(new_n16374), .O(new_n16377));
  inv1 g16184(.a(new_n16377), .O(new_n16378));
  nor2 g16185(.a(new_n16096), .b(new_n16092), .O(new_n16379));
  nor2 g16186(.a(new_n16379), .b(new_n16378), .O(new_n16380));
  inv1 g16187(.a(new_n16379), .O(new_n16381));
  nor2 g16188(.a(new_n16381), .b(new_n16377), .O(new_n16382));
  nor2 g16189(.a(new_n16382), .b(new_n16380), .O(new_n16383));
  inv1 g16190(.a(new_n16383), .O(\asquared[78] ));
  nor2 g16191(.a(new_n16370), .b(new_n16170), .O(new_n16385));
  nor2 g16192(.a(new_n16362), .b(new_n16272), .O(new_n16386));
  inv1 g16193(.a(new_n16386), .O(new_n16387));
  nor2 g16194(.a(new_n16247), .b(new_n16204), .O(new_n16388));
  nor2 g16195(.a(new_n16266), .b(new_n16260), .O(new_n16389));
  nor2 g16196(.a(new_n11596), .b(new_n800), .O(new_n16390));
  inv1 g16197(.a(new_n16390), .O(new_n16391));
  nor2 g16198(.a(new_n11186), .b(new_n847), .O(new_n16392));
  nor2 g16199(.a(new_n10895), .b(new_n941), .O(new_n16393));
  nor2 g16200(.a(new_n16393), .b(new_n16392), .O(new_n16394));
  nor2 g16201(.a(new_n11186), .b(new_n941), .O(new_n16395));
  inv1 g16202(.a(new_n16395), .O(new_n16396));
  nor2 g16203(.a(new_n16396), .b(new_n16108), .O(new_n16397));
  nor2 g16204(.a(new_n16397), .b(new_n16394), .O(new_n16398));
  nor2 g16205(.a(new_n16398), .b(new_n16391), .O(new_n16399));
  inv1 g16206(.a(new_n16398), .O(new_n16400));
  nor2 g16207(.a(new_n16400), .b(new_n16390), .O(new_n16401));
  nor2 g16208(.a(new_n16401), .b(new_n16399), .O(new_n16402));
  inv1 g16209(.a(new_n16402), .O(new_n16403));
  nor2 g16210(.a(new_n10320), .b(new_n1199), .O(new_n16404));
  nor2 g16211(.a(new_n16404), .b(new_n16338), .O(new_n16405));
  nor2 g16212(.a(new_n10320), .b(new_n1425), .O(new_n16406));
  inv1 g16213(.a(new_n16406), .O(new_n16407));
  nor2 g16214(.a(new_n16407), .b(new_n15838), .O(new_n16408));
  nor2 g16215(.a(new_n16408), .b(new_n16405), .O(new_n16409));
  inv1 g16216(.a(new_n16409), .O(new_n16410));
  nor2 g16217(.a(new_n16410), .b(new_n16182), .O(new_n16411));
  nor2 g16218(.a(new_n16409), .b(new_n16183), .O(new_n16412));
  nor2 g16219(.a(new_n16412), .b(new_n16411), .O(new_n16413));
  nor2 g16220(.a(new_n7537), .b(new_n2184), .O(new_n16414));
  inv1 g16221(.a(new_n16414), .O(new_n16415));
  nor2 g16222(.a(new_n7294), .b(new_n2433), .O(new_n16416));
  nor2 g16223(.a(new_n16416), .b(new_n16325), .O(new_n16417));
  inv1 g16224(.a(new_n16322), .O(new_n16418));
  nor2 g16225(.a(new_n7294), .b(new_n2506), .O(new_n16419));
  inv1 g16226(.a(new_n16419), .O(new_n16420));
  nor2 g16227(.a(new_n16420), .b(new_n16418), .O(new_n16421));
  nor2 g16228(.a(new_n16421), .b(new_n16417), .O(new_n16422));
  nor2 g16229(.a(new_n16422), .b(new_n16415), .O(new_n16423));
  inv1 g16230(.a(new_n16422), .O(new_n16424));
  nor2 g16231(.a(new_n16424), .b(new_n16414), .O(new_n16425));
  nor2 g16232(.a(new_n16425), .b(new_n16423), .O(new_n16426));
  nor2 g16233(.a(new_n16426), .b(new_n16413), .O(new_n16427));
  inv1 g16234(.a(new_n16413), .O(new_n16428));
  inv1 g16235(.a(new_n16426), .O(new_n16429));
  nor2 g16236(.a(new_n16429), .b(new_n16428), .O(new_n16430));
  nor2 g16237(.a(new_n16430), .b(new_n16427), .O(new_n16431));
  nor2 g16238(.a(new_n16431), .b(new_n16403), .O(new_n16432));
  inv1 g16239(.a(new_n16431), .O(new_n16433));
  nor2 g16240(.a(new_n16433), .b(new_n16402), .O(new_n16434));
  nor2 g16241(.a(new_n16434), .b(new_n16432), .O(new_n16435));
  inv1 g16242(.a(new_n16435), .O(new_n16436));
  nor2 g16243(.a(new_n8170), .b(new_n1903), .O(new_n16437));
  inv1 g16244(.a(new_n16437), .O(new_n16438));
  nor2 g16245(.a(new_n9156), .b(new_n1493), .O(new_n16439));
  nor2 g16246(.a(new_n16439), .b(new_n15030), .O(new_n16440));
  inv1 g16247(.a(new_n15811), .O(new_n16441));
  nor2 g16248(.a(new_n9156), .b(new_n1736), .O(new_n16442));
  inv1 g16249(.a(new_n16442), .O(new_n16443));
  nor2 g16250(.a(new_n16443), .b(new_n16441), .O(new_n16444));
  nor2 g16251(.a(new_n16444), .b(new_n16440), .O(new_n16445));
  nor2 g16252(.a(new_n16445), .b(new_n16438), .O(new_n16446));
  inv1 g16253(.a(new_n16445), .O(new_n16447));
  nor2 g16254(.a(new_n16447), .b(new_n16437), .O(new_n16448));
  nor2 g16255(.a(new_n16448), .b(new_n16446), .O(new_n16449));
  inv1 g16256(.a(new_n16449), .O(new_n16450));
  nor2 g16257(.a(new_n9873), .b(new_n1297), .O(new_n16451));
  nor2 g16258(.a(new_n6570), .b(new_n2826), .O(new_n16452));
  nor2 g16259(.a(new_n6893), .b(new_n2660), .O(new_n16453));
  nor2 g16260(.a(new_n16453), .b(new_n16452), .O(new_n16454));
  nor2 g16261(.a(new_n6893), .b(new_n2826), .O(new_n16455));
  inv1 g16262(.a(new_n16455), .O(new_n16456));
  nor2 g16263(.a(new_n16456), .b(new_n16002), .O(new_n16457));
  nor2 g16264(.a(new_n16457), .b(new_n16454), .O(new_n16458));
  inv1 g16265(.a(new_n16458), .O(new_n16459));
  nor2 g16266(.a(new_n16459), .b(new_n16451), .O(new_n16460));
  inv1 g16267(.a(new_n16451), .O(new_n16461));
  nor2 g16268(.a(new_n16458), .b(new_n16461), .O(new_n16462));
  nor2 g16269(.a(new_n16462), .b(new_n16460), .O(new_n16463));
  nor2 g16270(.a(new_n6274), .b(new_n3057), .O(new_n16464));
  nor2 g16271(.a(new_n5796), .b(new_n3533), .O(new_n16465));
  nor2 g16272(.a(new_n16465), .b(new_n16112), .O(new_n16466));
  inv1 g16273(.a(new_n16109), .O(new_n16467));
  nor2 g16274(.a(new_n5971), .b(new_n3533), .O(new_n16468));
  inv1 g16275(.a(new_n16468), .O(new_n16469));
  nor2 g16276(.a(new_n16469), .b(new_n16467), .O(new_n16470));
  nor2 g16277(.a(new_n16470), .b(new_n16466), .O(new_n16471));
  inv1 g16278(.a(new_n16471), .O(new_n16472));
  nor2 g16279(.a(new_n16472), .b(new_n16464), .O(new_n16473));
  inv1 g16280(.a(new_n16464), .O(new_n16474));
  nor2 g16281(.a(new_n16471), .b(new_n16474), .O(new_n16475));
  nor2 g16282(.a(new_n16475), .b(new_n16473), .O(new_n16476));
  nor2 g16283(.a(new_n16476), .b(new_n16463), .O(new_n16477));
  inv1 g16284(.a(new_n16463), .O(new_n16478));
  inv1 g16285(.a(new_n16476), .O(new_n16479));
  nor2 g16286(.a(new_n16479), .b(new_n16478), .O(new_n16480));
  nor2 g16287(.a(new_n16480), .b(new_n16477), .O(new_n16481));
  nor2 g16288(.a(new_n16481), .b(new_n16450), .O(new_n16482));
  inv1 g16289(.a(new_n16481), .O(new_n16483));
  nor2 g16290(.a(new_n16483), .b(new_n16449), .O(new_n16484));
  nor2 g16291(.a(new_n16484), .b(new_n16482), .O(new_n16485));
  inv1 g16292(.a(new_n16485), .O(new_n16486));
  nor2 g16293(.a(new_n16486), .b(new_n16436), .O(new_n16487));
  nor2 g16294(.a(new_n16485), .b(new_n16435), .O(new_n16488));
  nor2 g16295(.a(new_n16488), .b(new_n16487), .O(new_n16489));
  inv1 g16296(.a(new_n16489), .O(new_n16490));
  nor2 g16297(.a(new_n16490), .b(new_n16389), .O(new_n16491));
  inv1 g16298(.a(new_n16389), .O(new_n16492));
  nor2 g16299(.a(new_n16489), .b(new_n16492), .O(new_n16493));
  nor2 g16300(.a(new_n16493), .b(new_n16491), .O(new_n16494));
  inv1 g16301(.a(new_n16494), .O(new_n16495));
  nor2 g16302(.a(new_n16495), .b(new_n16388), .O(new_n16496));
  inv1 g16303(.a(new_n16388), .O(new_n16497));
  nor2 g16304(.a(new_n16494), .b(new_n16497), .O(new_n16498));
  nor2 g16305(.a(new_n16498), .b(new_n16496), .O(new_n16499));
  nor2 g16306(.a(new_n16499), .b(new_n16387), .O(new_n16500));
  inv1 g16307(.a(new_n16499), .O(new_n16501));
  nor2 g16308(.a(new_n16501), .b(new_n16386), .O(new_n16502));
  nor2 g16309(.a(new_n16502), .b(new_n16500), .O(new_n16503));
  inv1 g16310(.a(new_n16503), .O(new_n16504));
  nor2 g16311(.a(new_n16366), .b(new_n16252), .O(new_n16505));
  nor2 g16312(.a(new_n16505), .b(new_n16504), .O(new_n16506));
  inv1 g16313(.a(new_n16505), .O(new_n16507));
  nor2 g16314(.a(new_n16507), .b(new_n16503), .O(new_n16508));
  nor2 g16315(.a(new_n16508), .b(new_n16506), .O(new_n16509));
  inv1 g16316(.a(new_n16509), .O(new_n16510));
  nor2 g16317(.a(new_n16165), .b(new_n16160), .O(new_n16511));
  inv1 g16318(.a(new_n16511), .O(new_n16512));
  nor2 g16319(.a(new_n16353), .b(new_n16348), .O(new_n16513));
  inv1 g16320(.a(new_n16513), .O(new_n16514));
  nor2 g16321(.a(new_n16313), .b(new_n16300), .O(new_n16515));
  inv1 g16322(.a(new_n16515), .O(new_n16516));
  nor2 g16323(.a(new_n16516), .b(new_n16514), .O(new_n16517));
  nor2 g16324(.a(new_n16515), .b(new_n16513), .O(new_n16518));
  nor2 g16325(.a(new_n16518), .b(new_n16517), .O(new_n16519));
  nor2 g16326(.a(new_n16147), .b(new_n16142), .O(new_n16520));
  nor2 g16327(.a(new_n16520), .b(new_n16519), .O(new_n16521));
  inv1 g16328(.a(new_n16519), .O(new_n16522));
  inv1 g16329(.a(new_n16520), .O(new_n16523));
  nor2 g16330(.a(new_n16523), .b(new_n16522), .O(new_n16524));
  nor2 g16331(.a(new_n16524), .b(new_n16521), .O(new_n16525));
  inv1 g16332(.a(new_n16525), .O(new_n16526));
  nor2 g16333(.a(new_n16243), .b(new_n16240), .O(new_n16527));
  nor2 g16334(.a(new_n16527), .b(new_n16526), .O(new_n16528));
  inv1 g16335(.a(new_n16527), .O(new_n16529));
  nor2 g16336(.a(new_n16529), .b(new_n16525), .O(new_n16530));
  nor2 g16337(.a(new_n16530), .b(new_n16528), .O(new_n16531));
  inv1 g16338(.a(new_n16531), .O(new_n16532));
  nor2 g16339(.a(new_n16311), .b(new_n4425), .O(new_n16533));
  nor2 g16340(.a(new_n16287), .b(new_n16280), .O(new_n16534));
  nor2 g16341(.a(new_n16534), .b(new_n16533), .O(new_n16535));
  inv1 g16342(.a(new_n16533), .O(new_n16536));
  inv1 g16343(.a(new_n16534), .O(new_n16537));
  nor2 g16344(.a(new_n16537), .b(new_n16536), .O(new_n16538));
  nor2 g16345(.a(new_n16538), .b(new_n16535), .O(new_n16539));
  nor2 g16346(.a(new_n16126), .b(new_n16121), .O(new_n16540));
  nor2 g16347(.a(new_n16540), .b(new_n16539), .O(new_n16541));
  inv1 g16348(.a(new_n16539), .O(new_n16542));
  inv1 g16349(.a(new_n16540), .O(new_n16543));
  nor2 g16350(.a(new_n16543), .b(new_n16542), .O(new_n16544));
  nor2 g16351(.a(new_n16544), .b(new_n16541), .O(new_n16545));
  inv1 g16352(.a(new_n16545), .O(new_n16546));
  nor2 g16353(.a(new_n16298), .b(new_n16291), .O(new_n16547));
  nor2 g16354(.a(new_n16331), .b(new_n16324), .O(new_n16548));
  nor2 g16355(.a(new_n16548), .b(new_n16547), .O(new_n16549));
  inv1 g16356(.a(new_n16547), .O(new_n16550));
  inv1 g16357(.a(new_n16548), .O(new_n16551));
  nor2 g16358(.a(new_n16551), .b(new_n16550), .O(new_n16552));
  nor2 g16359(.a(new_n16552), .b(new_n16549), .O(new_n16553));
  nor2 g16360(.a(new_n16118), .b(new_n16110), .O(new_n16554));
  nor2 g16361(.a(new_n16554), .b(new_n16553), .O(new_n16555));
  inv1 g16362(.a(new_n16553), .O(new_n16556));
  inv1 g16363(.a(new_n16554), .O(new_n16557));
  nor2 g16364(.a(new_n16557), .b(new_n16556), .O(new_n16558));
  nor2 g16365(.a(new_n16558), .b(new_n16555), .O(new_n16559));
  nor2 g16366(.a(new_n16234), .b(new_n16228), .O(new_n16560));
  inv1 g16367(.a(new_n16560), .O(new_n16561));
  nor2 g16368(.a(new_n16561), .b(new_n16559), .O(new_n16562));
  inv1 g16369(.a(new_n16559), .O(new_n16563));
  nor2 g16370(.a(new_n16560), .b(new_n16563), .O(new_n16564));
  nor2 g16371(.a(new_n16564), .b(new_n16562), .O(new_n16565));
  inv1 g16372(.a(new_n16565), .O(new_n16566));
  nor2 g16373(.a(new_n16566), .b(new_n16546), .O(new_n16567));
  nor2 g16374(.a(new_n16565), .b(new_n16545), .O(new_n16568));
  nor2 g16375(.a(new_n16568), .b(new_n16567), .O(new_n16569));
  inv1 g16376(.a(new_n16569), .O(new_n16570));
  nor2 g16377(.a(new_n16570), .b(new_n16532), .O(new_n16571));
  nor2 g16378(.a(new_n16569), .b(new_n16531), .O(new_n16572));
  nor2 g16379(.a(new_n16572), .b(new_n16571), .O(new_n16573));
  nor2 g16380(.a(new_n16573), .b(new_n16512), .O(new_n16574));
  inv1 g16381(.a(new_n16573), .O(new_n16575));
  nor2 g16382(.a(new_n16575), .b(new_n16511), .O(new_n16576));
  nor2 g16383(.a(new_n16576), .b(new_n16574), .O(new_n16577));
  inv1 g16384(.a(new_n16577), .O(new_n16578));
  nor2 g16385(.a(new_n16220), .b(new_n16214), .O(new_n16579));
  inv1 g16386(.a(new_n16579), .O(new_n16580));
  nor2 g16387(.a(new_n8946), .b(new_n1647), .O(new_n16581));
  nor2 g16388(.a(new_n5393), .b(new_n3722), .O(new_n16582));
  nor2 g16389(.a(new_n5178), .b(new_n3870), .O(new_n16583));
  nor2 g16390(.a(new_n16583), .b(new_n16582), .O(new_n16584));
  nor2 g16391(.a(new_n5393), .b(new_n3870), .O(new_n16585));
  inv1 g16392(.a(new_n16585), .O(new_n16586));
  nor2 g16393(.a(new_n16586), .b(new_n16278), .O(new_n16587));
  nor2 g16394(.a(new_n16587), .b(new_n16584), .O(new_n16588));
  inv1 g16395(.a(new_n16588), .O(new_n16589));
  nor2 g16396(.a(new_n16589), .b(new_n16581), .O(new_n16590));
  inv1 g16397(.a(new_n16581), .O(new_n16591));
  nor2 g16398(.a(new_n16588), .b(new_n16591), .O(new_n16592));
  nor2 g16399(.a(new_n16592), .b(new_n16590), .O(new_n16593));
  nor2 g16400(.a(new_n8026), .b(new_n2121), .O(new_n16594));
  nor2 g16401(.a(new_n4682), .b(new_n4366), .O(new_n16595));
  nor2 g16402(.a(new_n16595), .b(new_n16594), .O(new_n16596));
  inv1 g16403(.a(new_n16594), .O(new_n16597));
  inv1 g16404(.a(new_n16595), .O(new_n16598));
  nor2 g16405(.a(new_n16598), .b(new_n16597), .O(new_n16599));
  nor2 g16406(.a(new_n16599), .b(new_n16596), .O(new_n16600));
  nor2 g16407(.a(new_n16600), .b(new_n16282), .O(new_n16601));
  inv1 g16408(.a(new_n16600), .O(new_n16602));
  nor2 g16409(.a(new_n16602), .b(new_n16281), .O(new_n16603));
  nor2 g16410(.a(new_n16603), .b(new_n16601), .O(new_n16604));
  nor2 g16411(.a(new_n16604), .b(new_n16593), .O(new_n16605));
  inv1 g16412(.a(new_n16593), .O(new_n16606));
  inv1 g16413(.a(new_n16604), .O(new_n16607));
  nor2 g16414(.a(new_n16607), .b(new_n16606), .O(new_n16608));
  nor2 g16415(.a(new_n16608), .b(new_n16605), .O(new_n16609));
  nor2 g16416(.a(new_n16609), .b(new_n16580), .O(new_n16610));
  inv1 g16417(.a(new_n16609), .O(new_n16611));
  nor2 g16418(.a(new_n16611), .b(new_n16579), .O(new_n16612));
  nor2 g16419(.a(new_n16612), .b(new_n16610), .O(new_n16613));
  inv1 g16420(.a(new_n16613), .O(new_n16614));
  nor2 g16421(.a(new_n16136), .b(new_n16133), .O(new_n16615));
  inv1 g16422(.a(new_n16615), .O(new_n16616));
  nor2 g16423(.a(new_n16344), .b(new_n16337), .O(new_n16617));
  nor2 g16424(.a(new_n16617), .b(new_n16616), .O(new_n16618));
  inv1 g16425(.a(new_n16617), .O(new_n16619));
  nor2 g16426(.a(new_n16619), .b(new_n16615), .O(new_n16620));
  nor2 g16427(.a(new_n16620), .b(new_n16618), .O(new_n16621));
  nor2 g16428(.a(new_n16189), .b(new_n16184), .O(new_n16622));
  inv1 g16429(.a(new_n16622), .O(new_n16623));
  nor2 g16430(.a(new_n16623), .b(new_n16621), .O(new_n16624));
  inv1 g16431(.a(new_n16621), .O(new_n16625));
  nor2 g16432(.a(new_n16622), .b(new_n16625), .O(new_n16626));
  nor2 g16433(.a(new_n16626), .b(new_n16624), .O(new_n16627));
  nor2 g16434(.a(new_n16200), .b(new_n16194), .O(new_n16628));
  inv1 g16435(.a(new_n16628), .O(new_n16629));
  nor2 g16436(.a(new_n16629), .b(new_n16627), .O(new_n16630));
  inv1 g16437(.a(new_n16627), .O(new_n16631));
  nor2 g16438(.a(new_n16628), .b(new_n16631), .O(new_n16632));
  nor2 g16439(.a(new_n16632), .b(new_n16630), .O(new_n16633));
  inv1 g16440(.a(new_n16633), .O(new_n16634));
  nor2 g16441(.a(new_n16634), .b(new_n16614), .O(new_n16635));
  nor2 g16442(.a(new_n16633), .b(new_n16613), .O(new_n16636));
  nor2 g16443(.a(new_n16636), .b(new_n16635), .O(new_n16637));
  inv1 g16444(.a(new_n16637), .O(new_n16638));
  nor2 g16445(.a(new_n16155), .b(new_n16149), .O(new_n16639));
  nor2 g16446(.a(new_n16358), .b(new_n16319), .O(new_n16640));
  nor2 g16447(.a(new_n16640), .b(new_n16639), .O(new_n16641));
  inv1 g16448(.a(new_n16639), .O(new_n16642));
  inv1 g16449(.a(new_n16640), .O(new_n16643));
  nor2 g16450(.a(new_n16643), .b(new_n16642), .O(new_n16644));
  nor2 g16451(.a(new_n16644), .b(new_n16641), .O(new_n16645));
  inv1 g16452(.a(new_n16645), .O(new_n16646));
  nor2 g16453(.a(new_n16646), .b(new_n16638), .O(new_n16647));
  nor2 g16454(.a(new_n16645), .b(new_n16637), .O(new_n16648));
  nor2 g16455(.a(new_n16648), .b(new_n16647), .O(new_n16649));
  inv1 g16456(.a(new_n16649), .O(new_n16650));
  nor2 g16457(.a(new_n16650), .b(new_n16578), .O(new_n16651));
  nor2 g16458(.a(new_n16649), .b(new_n16577), .O(new_n16652));
  nor2 g16459(.a(new_n16652), .b(new_n16651), .O(new_n16653));
  inv1 g16460(.a(new_n16653), .O(new_n16654));
  nor2 g16461(.a(new_n16654), .b(new_n16510), .O(new_n16655));
  nor2 g16462(.a(new_n16653), .b(new_n16509), .O(new_n16656));
  nor2 g16463(.a(new_n16656), .b(new_n16655), .O(new_n16657));
  inv1 g16464(.a(new_n16657), .O(new_n16658));
  nor2 g16465(.a(new_n16658), .b(new_n16385), .O(new_n16659));
  inv1 g16466(.a(new_n16385), .O(new_n16660));
  nor2 g16467(.a(new_n16657), .b(new_n16660), .O(new_n16661));
  nor2 g16468(.a(new_n16661), .b(new_n16659), .O(new_n16662));
  inv1 g16469(.a(new_n16662), .O(new_n16663));
  nor2 g16470(.a(new_n16380), .b(new_n16376), .O(new_n16664));
  nor2 g16471(.a(new_n16664), .b(new_n16663), .O(new_n16665));
  inv1 g16472(.a(new_n16664), .O(new_n16666));
  nor2 g16473(.a(new_n16666), .b(new_n16662), .O(new_n16667));
  nor2 g16474(.a(new_n16667), .b(new_n16665), .O(new_n16668));
  inv1 g16475(.a(new_n16668), .O(\asquared[79] ));
  nor2 g16476(.a(new_n16655), .b(new_n16506), .O(new_n16670));
  nor2 g16477(.a(new_n16647), .b(new_n16641), .O(new_n16671));
  inv1 g16478(.a(new_n16671), .O(new_n16672));
  nor2 g16479(.a(new_n16491), .b(new_n16487), .O(new_n16673));
  inv1 g16480(.a(new_n16673), .O(new_n16674));
  nor2 g16481(.a(new_n16425), .b(new_n16417), .O(new_n16675));
  nor2 g16482(.a(new_n16411), .b(new_n16405), .O(new_n16676));
  nor2 g16483(.a(new_n16676), .b(new_n16675), .O(new_n16677));
  inv1 g16484(.a(new_n16675), .O(new_n16678));
  inv1 g16485(.a(new_n16676), .O(new_n16679));
  nor2 g16486(.a(new_n16679), .b(new_n16678), .O(new_n16680));
  nor2 g16487(.a(new_n16680), .b(new_n16677), .O(new_n16681));
  nor2 g16488(.a(new_n16448), .b(new_n16440), .O(new_n16682));
  nor2 g16489(.a(new_n16682), .b(new_n16681), .O(new_n16683));
  inv1 g16490(.a(new_n16681), .O(new_n16684));
  inv1 g16491(.a(new_n16682), .O(new_n16685));
  nor2 g16492(.a(new_n16685), .b(new_n16684), .O(new_n16686));
  nor2 g16493(.a(new_n16686), .b(new_n16683), .O(new_n16687));
  nor2 g16494(.a(new_n16612), .b(new_n16605), .O(new_n16688));
  inv1 g16495(.a(new_n16688), .O(new_n16689));
  nor2 g16496(.a(new_n16689), .b(new_n16687), .O(new_n16690));
  inv1 g16497(.a(new_n16687), .O(new_n16691));
  nor2 g16498(.a(new_n16688), .b(new_n16691), .O(new_n16692));
  nor2 g16499(.a(new_n16692), .b(new_n16690), .O(new_n16693));
  inv1 g16500(.a(new_n16693), .O(new_n16694));
  nor2 g16501(.a(new_n16626), .b(new_n16620), .O(new_n16695));
  inv1 g16502(.a(new_n16695), .O(new_n16696));
  nor2 g16503(.a(new_n11596), .b(new_n847), .O(new_n16697));
  nor2 g16504(.a(new_n5796), .b(new_n3722), .O(new_n16698));
  nor2 g16505(.a(new_n16698), .b(new_n16468), .O(new_n16699));
  inv1 g16506(.a(new_n16465), .O(new_n16700));
  nor2 g16507(.a(new_n5971), .b(new_n3722), .O(new_n16701));
  inv1 g16508(.a(new_n16701), .O(new_n16702));
  nor2 g16509(.a(new_n16702), .b(new_n16700), .O(new_n16703));
  nor2 g16510(.a(new_n16703), .b(new_n16699), .O(new_n16704));
  inv1 g16511(.a(new_n16704), .O(new_n16705));
  nor2 g16512(.a(new_n16705), .b(new_n16697), .O(new_n16706));
  inv1 g16513(.a(new_n16697), .O(new_n16707));
  nor2 g16514(.a(new_n16704), .b(new_n16707), .O(new_n16708));
  nor2 g16515(.a(new_n16708), .b(new_n16706), .O(new_n16709));
  nor2 g16516(.a(new_n9156), .b(new_n1647), .O(new_n16710));
  nor2 g16517(.a(new_n8026), .b(new_n2184), .O(new_n16711));
  nor2 g16518(.a(new_n16711), .b(new_n16710), .O(new_n16712));
  nor2 g16519(.a(new_n9156), .b(new_n2184), .O(new_n16713));
  inv1 g16520(.a(new_n16713), .O(new_n16714));
  nor2 g16521(.a(new_n16714), .b(new_n15616), .O(new_n16715));
  nor2 g16522(.a(new_n16715), .b(new_n16712), .O(new_n16716));
  nor2 g16523(.a(new_n16716), .b(new_n16586), .O(new_n16717));
  inv1 g16524(.a(new_n16716), .O(new_n16718));
  nor2 g16525(.a(new_n16718), .b(new_n16585), .O(new_n16719));
  nor2 g16526(.a(new_n16719), .b(new_n16717), .O(new_n16720));
  nor2 g16527(.a(new_n16720), .b(new_n16709), .O(new_n16721));
  inv1 g16528(.a(new_n16709), .O(new_n16722));
  inv1 g16529(.a(new_n16720), .O(new_n16723));
  nor2 g16530(.a(new_n16723), .b(new_n16722), .O(new_n16724));
  nor2 g16531(.a(new_n16724), .b(new_n16721), .O(new_n16725));
  nor2 g16532(.a(new_n16725), .b(new_n16696), .O(new_n16726));
  inv1 g16533(.a(new_n16725), .O(new_n16727));
  nor2 g16534(.a(new_n16727), .b(new_n16695), .O(new_n16728));
  nor2 g16535(.a(new_n16728), .b(new_n16726), .O(new_n16729));
  inv1 g16536(.a(new_n16729), .O(new_n16730));
  nor2 g16537(.a(new_n16730), .b(new_n16694), .O(new_n16731));
  nor2 g16538(.a(new_n16729), .b(new_n16693), .O(new_n16732));
  nor2 g16539(.a(new_n16732), .b(new_n16731), .O(new_n16733));
  nor2 g16540(.a(new_n16733), .b(new_n16674), .O(new_n16734));
  inv1 g16541(.a(new_n16733), .O(new_n16735));
  nor2 g16542(.a(new_n16735), .b(new_n16673), .O(new_n16736));
  nor2 g16543(.a(new_n16736), .b(new_n16734), .O(new_n16737));
  inv1 g16544(.a(new_n16737), .O(new_n16738));
  nor2 g16545(.a(new_n10895), .b(new_n1086), .O(new_n16739));
  inv1 g16546(.a(new_n16739), .O(new_n16740));
  nor2 g16547(.a(new_n16603), .b(new_n16596), .O(new_n16741));
  inv1 g16548(.a(new_n16741), .O(new_n16742));
  nor2 g16549(.a(new_n16742), .b(new_n16740), .O(new_n16743));
  nor2 g16550(.a(new_n16741), .b(new_n16739), .O(new_n16744));
  nor2 g16551(.a(new_n16744), .b(new_n16743), .O(new_n16745));
  nor2 g16552(.a(new_n16590), .b(new_n16584), .O(new_n16746));
  nor2 g16553(.a(new_n16746), .b(new_n16745), .O(new_n16747));
  inv1 g16554(.a(new_n16745), .O(new_n16748));
  inv1 g16555(.a(new_n16746), .O(new_n16749));
  nor2 g16556(.a(new_n16749), .b(new_n16748), .O(new_n16750));
  nor2 g16557(.a(new_n16750), .b(new_n16747), .O(new_n16751));
  inv1 g16558(.a(new_n16751), .O(new_n16752));
  nor2 g16559(.a(new_n16401), .b(new_n16394), .O(new_n16753));
  nor2 g16560(.a(new_n16460), .b(new_n16454), .O(new_n16754));
  nor2 g16561(.a(new_n16754), .b(new_n16753), .O(new_n16755));
  inv1 g16562(.a(new_n16753), .O(new_n16756));
  inv1 g16563(.a(new_n16754), .O(new_n16757));
  nor2 g16564(.a(new_n16757), .b(new_n16756), .O(new_n16758));
  nor2 g16565(.a(new_n16758), .b(new_n16755), .O(new_n16759));
  nor2 g16566(.a(new_n16473), .b(new_n16466), .O(new_n16760));
  nor2 g16567(.a(new_n16760), .b(new_n16759), .O(new_n16761));
  inv1 g16568(.a(new_n16759), .O(new_n16762));
  inv1 g16569(.a(new_n16760), .O(new_n16763));
  nor2 g16570(.a(new_n16763), .b(new_n16762), .O(new_n16764));
  nor2 g16571(.a(new_n16764), .b(new_n16761), .O(new_n16765));
  inv1 g16572(.a(new_n16765), .O(new_n16766));
  nor2 g16573(.a(new_n16766), .b(new_n16752), .O(new_n16767));
  nor2 g16574(.a(new_n16765), .b(new_n16751), .O(new_n16768));
  nor2 g16575(.a(new_n16768), .b(new_n16767), .O(new_n16769));
  inv1 g16576(.a(new_n16769), .O(new_n16770));
  nor2 g16577(.a(new_n16484), .b(new_n16477), .O(new_n16771));
  nor2 g16578(.a(new_n16771), .b(new_n16770), .O(new_n16772));
  inv1 g16579(.a(new_n16771), .O(new_n16773));
  nor2 g16580(.a(new_n16773), .b(new_n16769), .O(new_n16774));
  nor2 g16581(.a(new_n16774), .b(new_n16772), .O(new_n16775));
  inv1 g16582(.a(new_n16775), .O(new_n16776));
  nor2 g16583(.a(new_n16776), .b(new_n16738), .O(new_n16777));
  nor2 g16584(.a(new_n16775), .b(new_n16737), .O(new_n16778));
  nor2 g16585(.a(new_n16778), .b(new_n16777), .O(new_n16779));
  nor2 g16586(.a(new_n16779), .b(new_n16672), .O(new_n16780));
  inv1 g16587(.a(new_n16779), .O(new_n16781));
  nor2 g16588(.a(new_n16781), .b(new_n16671), .O(new_n16782));
  nor2 g16589(.a(new_n16782), .b(new_n16780), .O(new_n16783));
  nor2 g16590(.a(new_n16502), .b(new_n16496), .O(new_n16784));
  inv1 g16591(.a(new_n16784), .O(new_n16785));
  nor2 g16592(.a(new_n16785), .b(new_n16783), .O(new_n16786));
  inv1 g16593(.a(new_n16783), .O(new_n16787));
  nor2 g16594(.a(new_n16784), .b(new_n16787), .O(new_n16788));
  nor2 g16595(.a(new_n16788), .b(new_n16786), .O(new_n16789));
  inv1 g16596(.a(new_n16789), .O(new_n16790));
  nor2 g16597(.a(new_n16571), .b(new_n16528), .O(new_n16791));
  inv1 g16598(.a(new_n16791), .O(new_n16792));
  nor2 g16599(.a(new_n16567), .b(new_n16564), .O(new_n16793));
  nor2 g16600(.a(new_n7537), .b(new_n2433), .O(new_n16794));
  inv1 g16601(.a(new_n16794), .O(new_n16795));
  nor2 g16602(.a(new_n11186), .b(new_n4682), .O(new_n16796));
  inv1 g16603(.a(new_n16796), .O(new_n16797));
  nor2 g16604(.a(new_n16797), .b(new_n941), .O(new_n16798));
  nor2 g16605(.a(new_n16395), .b(\a[40] ), .O(new_n16799));
  nor2 g16606(.a(new_n16799), .b(new_n16795), .O(new_n16800));
  inv1 g16607(.a(new_n16800), .O(new_n16801));
  nor2 g16608(.a(new_n16801), .b(new_n16798), .O(new_n16802));
  nor2 g16609(.a(new_n16802), .b(new_n16795), .O(new_n16803));
  nor2 g16610(.a(new_n16800), .b(new_n16798), .O(new_n16804));
  inv1 g16611(.a(new_n16804), .O(new_n16805));
  nor2 g16612(.a(new_n16805), .b(new_n16799), .O(new_n16806));
  nor2 g16613(.a(new_n16806), .b(new_n16803), .O(new_n16807));
  nor2 g16614(.a(new_n8946), .b(new_n1736), .O(new_n16808));
  nor2 g16615(.a(new_n8170), .b(new_n2121), .O(new_n16809));
  nor2 g16616(.a(new_n8476), .b(new_n1903), .O(new_n16810));
  nor2 g16617(.a(new_n16810), .b(new_n16809), .O(new_n16811));
  nor2 g16618(.a(new_n8476), .b(new_n2121), .O(new_n16812));
  inv1 g16619(.a(new_n16812), .O(new_n16813));
  nor2 g16620(.a(new_n16813), .b(new_n16438), .O(new_n16814));
  nor2 g16621(.a(new_n16814), .b(new_n16811), .O(new_n16815));
  inv1 g16622(.a(new_n16815), .O(new_n16816));
  nor2 g16623(.a(new_n16816), .b(new_n16808), .O(new_n16817));
  inv1 g16624(.a(new_n16808), .O(new_n16818));
  nor2 g16625(.a(new_n16815), .b(new_n16818), .O(new_n16819));
  nor2 g16626(.a(new_n16819), .b(new_n16817), .O(new_n16820));
  nor2 g16627(.a(new_n5178), .b(new_n4093), .O(new_n16821));
  inv1 g16628(.a(new_n16821), .O(new_n16822));
  nor2 g16629(.a(new_n4954), .b(new_n4366), .O(new_n16823));
  nor2 g16630(.a(new_n4682), .b(new_n4425), .O(new_n16824));
  nor2 g16631(.a(new_n16824), .b(new_n16823), .O(new_n16825));
  nor2 g16632(.a(new_n4954), .b(new_n4425), .O(new_n16826));
  inv1 g16633(.a(new_n16826), .O(new_n16827));
  nor2 g16634(.a(new_n16827), .b(new_n16598), .O(new_n16828));
  nor2 g16635(.a(new_n16828), .b(new_n16825), .O(new_n16829));
  nor2 g16636(.a(new_n16829), .b(new_n16822), .O(new_n16830));
  inv1 g16637(.a(new_n16829), .O(new_n16831));
  nor2 g16638(.a(new_n16831), .b(new_n16821), .O(new_n16832));
  nor2 g16639(.a(new_n16832), .b(new_n16830), .O(new_n16833));
  nor2 g16640(.a(new_n16833), .b(new_n16820), .O(new_n16834));
  inv1 g16641(.a(new_n16820), .O(new_n16835));
  inv1 g16642(.a(new_n16833), .O(new_n16836));
  nor2 g16643(.a(new_n16836), .b(new_n16835), .O(new_n16837));
  nor2 g16644(.a(new_n16837), .b(new_n16834), .O(new_n16838));
  inv1 g16645(.a(new_n16838), .O(new_n16839));
  nor2 g16646(.a(new_n16839), .b(new_n16807), .O(new_n16840));
  inv1 g16647(.a(new_n16807), .O(new_n16841));
  nor2 g16648(.a(new_n16838), .b(new_n16841), .O(new_n16842));
  nor2 g16649(.a(new_n16842), .b(new_n16840), .O(new_n16843));
  nor2 g16650(.a(new_n6274), .b(new_n3231), .O(new_n16844));
  nor2 g16651(.a(new_n6570), .b(new_n3057), .O(new_n16845));
  nor2 g16652(.a(new_n16845), .b(new_n16844), .O(new_n16846));
  nor2 g16653(.a(new_n6570), .b(new_n3231), .O(new_n16847));
  inv1 g16654(.a(new_n16847), .O(new_n16848));
  nor2 g16655(.a(new_n16848), .b(new_n16474), .O(new_n16849));
  nor2 g16656(.a(new_n16849), .b(new_n16846), .O(new_n16850));
  nor2 g16657(.a(new_n16850), .b(new_n16456), .O(new_n16851));
  inv1 g16658(.a(new_n16850), .O(new_n16852));
  nor2 g16659(.a(new_n16852), .b(new_n16455), .O(new_n16853));
  nor2 g16660(.a(new_n16853), .b(new_n16851), .O(new_n16854));
  inv1 g16661(.a(new_n16854), .O(new_n16855));
  nor2 g16662(.a(new_n10468), .b(new_n1199), .O(new_n16856));
  nor2 g16663(.a(new_n10320), .b(new_n1297), .O(new_n16857));
  nor2 g16664(.a(new_n9873), .b(new_n1425), .O(new_n16858));
  nor2 g16665(.a(new_n16858), .b(new_n16857), .O(new_n16859));
  nor2 g16666(.a(new_n16461), .b(new_n16407), .O(new_n16860));
  nor2 g16667(.a(new_n16860), .b(new_n16859), .O(new_n16861));
  inv1 g16668(.a(new_n16861), .O(new_n16862));
  nor2 g16669(.a(new_n16862), .b(new_n16856), .O(new_n16863));
  inv1 g16670(.a(new_n16856), .O(new_n16864));
  nor2 g16671(.a(new_n16861), .b(new_n16864), .O(new_n16865));
  nor2 g16672(.a(new_n16865), .b(new_n16863), .O(new_n16866));
  nor2 g16673(.a(new_n9658), .b(new_n1493), .O(new_n16867));
  inv1 g16674(.a(new_n16867), .O(new_n16868));
  nor2 g16675(.a(new_n6958), .b(new_n2660), .O(new_n16869));
  nor2 g16676(.a(new_n16869), .b(new_n16419), .O(new_n16870));
  nor2 g16677(.a(new_n7294), .b(new_n2660), .O(new_n16871));
  inv1 g16678(.a(new_n16871), .O(new_n16872));
  nor2 g16679(.a(new_n16872), .b(new_n16326), .O(new_n16873));
  nor2 g16680(.a(new_n16873), .b(new_n16870), .O(new_n16874));
  nor2 g16681(.a(new_n16874), .b(new_n16868), .O(new_n16875));
  inv1 g16682(.a(new_n16874), .O(new_n16876));
  nor2 g16683(.a(new_n16876), .b(new_n16867), .O(new_n16877));
  nor2 g16684(.a(new_n16877), .b(new_n16875), .O(new_n16878));
  nor2 g16685(.a(new_n16878), .b(new_n16866), .O(new_n16879));
  inv1 g16686(.a(new_n16866), .O(new_n16880));
  inv1 g16687(.a(new_n16878), .O(new_n16881));
  nor2 g16688(.a(new_n16881), .b(new_n16880), .O(new_n16882));
  nor2 g16689(.a(new_n16882), .b(new_n16879), .O(new_n16883));
  nor2 g16690(.a(new_n16883), .b(new_n16855), .O(new_n16884));
  inv1 g16691(.a(new_n16883), .O(new_n16885));
  nor2 g16692(.a(new_n16885), .b(new_n16854), .O(new_n16886));
  nor2 g16693(.a(new_n16886), .b(new_n16884), .O(new_n16887));
  nor2 g16694(.a(new_n16887), .b(new_n16843), .O(new_n16888));
  inv1 g16695(.a(new_n16843), .O(new_n16889));
  inv1 g16696(.a(new_n16887), .O(new_n16890));
  nor2 g16697(.a(new_n16890), .b(new_n16889), .O(new_n16891));
  nor2 g16698(.a(new_n16891), .b(new_n16888), .O(new_n16892));
  inv1 g16699(.a(new_n16892), .O(new_n16893));
  nor2 g16700(.a(new_n16893), .b(new_n16793), .O(new_n16894));
  inv1 g16701(.a(new_n16793), .O(new_n16895));
  nor2 g16702(.a(new_n16892), .b(new_n16895), .O(new_n16896));
  nor2 g16703(.a(new_n16896), .b(new_n16894), .O(new_n16897));
  nor2 g16704(.a(new_n16897), .b(new_n16792), .O(new_n16898));
  inv1 g16705(.a(new_n16897), .O(new_n16899));
  nor2 g16706(.a(new_n16899), .b(new_n16791), .O(new_n16900));
  nor2 g16707(.a(new_n16900), .b(new_n16898), .O(new_n16901));
  inv1 g16708(.a(new_n16901), .O(new_n16902));
  nor2 g16709(.a(new_n16558), .b(new_n16552), .O(new_n16903));
  inv1 g16710(.a(new_n16903), .O(new_n16904));
  nor2 g16711(.a(new_n16544), .b(new_n16538), .O(new_n16905));
  inv1 g16712(.a(new_n16905), .O(new_n16906));
  nor2 g16713(.a(new_n16906), .b(new_n16904), .O(new_n16907));
  nor2 g16714(.a(new_n16905), .b(new_n16903), .O(new_n16908));
  nor2 g16715(.a(new_n16908), .b(new_n16907), .O(new_n16909));
  nor2 g16716(.a(new_n16434), .b(new_n16427), .O(new_n16910));
  inv1 g16717(.a(new_n16910), .O(new_n16911));
  nor2 g16718(.a(new_n16911), .b(new_n16909), .O(new_n16912));
  inv1 g16719(.a(new_n16909), .O(new_n16913));
  nor2 g16720(.a(new_n16910), .b(new_n16913), .O(new_n16914));
  nor2 g16721(.a(new_n16914), .b(new_n16912), .O(new_n16915));
  nor2 g16722(.a(new_n16524), .b(new_n16518), .O(new_n16916));
  inv1 g16723(.a(new_n16916), .O(new_n16917));
  nor2 g16724(.a(new_n16917), .b(new_n16915), .O(new_n16918));
  inv1 g16725(.a(new_n16915), .O(new_n16919));
  nor2 g16726(.a(new_n16916), .b(new_n16919), .O(new_n16920));
  nor2 g16727(.a(new_n16920), .b(new_n16918), .O(new_n16921));
  inv1 g16728(.a(new_n16921), .O(new_n16922));
  nor2 g16729(.a(new_n16635), .b(new_n16632), .O(new_n16923));
  nor2 g16730(.a(new_n16923), .b(new_n16922), .O(new_n16924));
  inv1 g16731(.a(new_n16923), .O(new_n16925));
  nor2 g16732(.a(new_n16925), .b(new_n16921), .O(new_n16926));
  nor2 g16733(.a(new_n16926), .b(new_n16924), .O(new_n16927));
  inv1 g16734(.a(new_n16927), .O(new_n16928));
  nor2 g16735(.a(new_n16928), .b(new_n16902), .O(new_n16929));
  nor2 g16736(.a(new_n16927), .b(new_n16901), .O(new_n16930));
  nor2 g16737(.a(new_n16930), .b(new_n16929), .O(new_n16931));
  inv1 g16738(.a(new_n16931), .O(new_n16932));
  nor2 g16739(.a(new_n16651), .b(new_n16576), .O(new_n16933));
  nor2 g16740(.a(new_n16933), .b(new_n16932), .O(new_n16934));
  inv1 g16741(.a(new_n16933), .O(new_n16935));
  nor2 g16742(.a(new_n16935), .b(new_n16931), .O(new_n16936));
  nor2 g16743(.a(new_n16936), .b(new_n16934), .O(new_n16937));
  inv1 g16744(.a(new_n16937), .O(new_n16938));
  nor2 g16745(.a(new_n16938), .b(new_n16790), .O(new_n16939));
  nor2 g16746(.a(new_n16937), .b(new_n16789), .O(new_n16940));
  nor2 g16747(.a(new_n16940), .b(new_n16939), .O(new_n16941));
  inv1 g16748(.a(new_n16941), .O(new_n16942));
  nor2 g16749(.a(new_n16942), .b(new_n16670), .O(new_n16943));
  inv1 g16750(.a(new_n16670), .O(new_n16944));
  nor2 g16751(.a(new_n16941), .b(new_n16944), .O(new_n16945));
  nor2 g16752(.a(new_n16945), .b(new_n16943), .O(new_n16946));
  inv1 g16753(.a(new_n16946), .O(new_n16947));
  nor2 g16754(.a(new_n16665), .b(new_n16661), .O(new_n16948));
  nor2 g16755(.a(new_n16948), .b(new_n16947), .O(new_n16949));
  inv1 g16756(.a(new_n16948), .O(new_n16950));
  nor2 g16757(.a(new_n16950), .b(new_n16946), .O(new_n16951));
  nor2 g16758(.a(new_n16951), .b(new_n16949), .O(new_n16952));
  inv1 g16759(.a(new_n16952), .O(\asquared[80] ));
  nor2 g16760(.a(new_n16939), .b(new_n16934), .O(new_n16954));
  inv1 g16761(.a(new_n16954), .O(new_n16955));
  nor2 g16762(.a(new_n16788), .b(new_n16782), .O(new_n16956));
  inv1 g16763(.a(new_n16956), .O(new_n16957));
  nor2 g16764(.a(new_n16777), .b(new_n16736), .O(new_n16958));
  nor2 g16765(.a(new_n16924), .b(new_n16920), .O(new_n16959));
  nor2 g16766(.a(new_n10895), .b(new_n1199), .O(new_n16960));
  nor2 g16767(.a(new_n11186), .b(new_n1086), .O(new_n16961));
  nor2 g16768(.a(new_n16961), .b(new_n16960), .O(new_n16962));
  nor2 g16769(.a(new_n11186), .b(new_n1199), .O(new_n16963));
  inv1 g16770(.a(new_n16963), .O(new_n16964));
  nor2 g16771(.a(new_n16964), .b(new_n16740), .O(new_n16965));
  nor2 g16772(.a(new_n16965), .b(new_n16962), .O(new_n16966));
  inv1 g16773(.a(new_n16966), .O(new_n16967));
  nor2 g16774(.a(new_n16967), .b(new_n16804), .O(new_n16968));
  nor2 g16775(.a(new_n16966), .b(new_n16805), .O(new_n16969));
  nor2 g16776(.a(new_n16969), .b(new_n16968), .O(new_n16970));
  inv1 g16777(.a(new_n16970), .O(new_n16971));
  nor2 g16778(.a(new_n11596), .b(new_n941), .O(new_n16972));
  nor2 g16779(.a(new_n7537), .b(new_n2506), .O(new_n16973));
  nor2 g16780(.a(new_n16973), .b(new_n16972), .O(new_n16974));
  nor2 g16781(.a(new_n11596), .b(new_n2506), .O(new_n16975));
  inv1 g16782(.a(new_n16975), .O(new_n16976));
  nor2 g16783(.a(new_n16976), .b(new_n9506), .O(new_n16977));
  nor2 g16784(.a(new_n16977), .b(new_n16974), .O(new_n16978));
  inv1 g16785(.a(new_n16978), .O(new_n16979));
  nor2 g16786(.a(new_n16979), .b(new_n16847), .O(new_n16980));
  nor2 g16787(.a(new_n16978), .b(new_n16848), .O(new_n16981));
  nor2 g16788(.a(new_n16981), .b(new_n16980), .O(new_n16982));
  nor2 g16789(.a(new_n6274), .b(new_n3533), .O(new_n16983));
  inv1 g16790(.a(new_n16983), .O(new_n16984));
  nor2 g16791(.a(new_n5796), .b(new_n3870), .O(new_n16985));
  nor2 g16792(.a(new_n16985), .b(new_n16701), .O(new_n16986));
  inv1 g16793(.a(new_n16698), .O(new_n16987));
  nor2 g16794(.a(new_n5971), .b(new_n3870), .O(new_n16988));
  inv1 g16795(.a(new_n16988), .O(new_n16989));
  nor2 g16796(.a(new_n16989), .b(new_n16987), .O(new_n16990));
  nor2 g16797(.a(new_n16990), .b(new_n16986), .O(new_n16991));
  nor2 g16798(.a(new_n16991), .b(new_n16984), .O(new_n16992));
  inv1 g16799(.a(new_n16991), .O(new_n16993));
  nor2 g16800(.a(new_n16993), .b(new_n16983), .O(new_n16994));
  nor2 g16801(.a(new_n16994), .b(new_n16992), .O(new_n16995));
  nor2 g16802(.a(new_n16995), .b(new_n16982), .O(new_n16996));
  inv1 g16803(.a(new_n16982), .O(new_n16997));
  inv1 g16804(.a(new_n16995), .O(new_n16998));
  nor2 g16805(.a(new_n16998), .b(new_n16997), .O(new_n16999));
  nor2 g16806(.a(new_n16999), .b(new_n16996), .O(new_n17000));
  inv1 g16807(.a(new_n17000), .O(new_n17001));
  nor2 g16808(.a(new_n17001), .b(new_n16971), .O(new_n17002));
  nor2 g16809(.a(new_n17000), .b(new_n16970), .O(new_n17003));
  nor2 g16810(.a(new_n17003), .b(new_n17002), .O(new_n17004));
  inv1 g16811(.a(new_n17004), .O(new_n17005));
  nor2 g16812(.a(new_n9873), .b(new_n1493), .O(new_n17006));
  nor2 g16813(.a(new_n17006), .b(new_n16406), .O(new_n17007));
  inv1 g16814(.a(new_n16858), .O(new_n17008));
  nor2 g16815(.a(new_n10320), .b(new_n1493), .O(new_n17009));
  inv1 g16816(.a(new_n17009), .O(new_n17010));
  nor2 g16817(.a(new_n17010), .b(new_n17008), .O(new_n17011));
  nor2 g16818(.a(new_n17011), .b(new_n17007), .O(new_n17012));
  nor2 g16819(.a(new_n10468), .b(new_n1297), .O(new_n17013));
  nor2 g16820(.a(new_n17013), .b(new_n17012), .O(new_n17014));
  inv1 g16821(.a(new_n17012), .O(new_n17015));
  inv1 g16822(.a(new_n17013), .O(new_n17016));
  nor2 g16823(.a(new_n17016), .b(new_n17015), .O(new_n17017));
  nor2 g16824(.a(new_n17017), .b(new_n17014), .O(new_n17018));
  inv1 g16825(.a(new_n17018), .O(new_n17019));
  nor2 g16826(.a(new_n16832), .b(new_n16825), .O(new_n17020));
  inv1 g16827(.a(new_n17020), .O(new_n17021));
  nor2 g16828(.a(new_n17021), .b(new_n17019), .O(new_n17022));
  nor2 g16829(.a(new_n17020), .b(new_n17018), .O(new_n17023));
  nor2 g16830(.a(new_n17023), .b(new_n17022), .O(new_n17024));
  inv1 g16831(.a(new_n17024), .O(new_n17025));
  nor2 g16832(.a(new_n6958), .b(new_n2826), .O(new_n17026));
  nor2 g16833(.a(new_n6893), .b(new_n3057), .O(new_n17027));
  nor2 g16834(.a(new_n17027), .b(new_n17026), .O(new_n17028));
  nor2 g16835(.a(new_n6958), .b(new_n3057), .O(new_n17029));
  inv1 g16836(.a(new_n17029), .O(new_n17030));
  nor2 g16837(.a(new_n17030), .b(new_n16456), .O(new_n17031));
  nor2 g16838(.a(new_n17031), .b(new_n17028), .O(new_n17032));
  nor2 g16839(.a(new_n17032), .b(new_n16872), .O(new_n17033));
  inv1 g16840(.a(new_n17032), .O(new_n17034));
  nor2 g16841(.a(new_n17034), .b(new_n16871), .O(new_n17035));
  nor2 g16842(.a(new_n17035), .b(new_n17033), .O(new_n17036));
  nor2 g16843(.a(new_n17036), .b(new_n17025), .O(new_n17037));
  inv1 g16844(.a(new_n17036), .O(new_n17038));
  nor2 g16845(.a(new_n17038), .b(new_n17024), .O(new_n17039));
  nor2 g16846(.a(new_n17039), .b(new_n17037), .O(new_n17040));
  inv1 g16847(.a(new_n17040), .O(new_n17041));
  nor2 g16848(.a(new_n8170), .b(new_n2184), .O(new_n17042));
  nor2 g16849(.a(new_n8026), .b(new_n2433), .O(new_n17043));
  nor2 g16850(.a(new_n17043), .b(new_n17042), .O(new_n17044));
  inv1 g16851(.a(new_n16711), .O(new_n17045));
  nor2 g16852(.a(new_n8170), .b(new_n2433), .O(new_n17046));
  inv1 g16853(.a(new_n17046), .O(new_n17047));
  nor2 g16854(.a(new_n17047), .b(new_n17045), .O(new_n17048));
  nor2 g16855(.a(new_n17048), .b(new_n17044), .O(new_n17049));
  nor2 g16856(.a(new_n17049), .b(new_n16827), .O(new_n17050));
  inv1 g16857(.a(new_n17049), .O(new_n17051));
  nor2 g16858(.a(new_n17051), .b(new_n16826), .O(new_n17052));
  nor2 g16859(.a(new_n17052), .b(new_n17050), .O(new_n17053));
  inv1 g16860(.a(new_n17053), .O(new_n17054));
  nor2 g16861(.a(new_n9658), .b(new_n1647), .O(new_n17055));
  nor2 g16862(.a(new_n16812), .b(new_n16442), .O(new_n17056));
  nor2 g16863(.a(new_n9156), .b(new_n2121), .O(new_n17057));
  inv1 g16864(.a(new_n17057), .O(new_n17058));
  nor2 g16865(.a(new_n17058), .b(new_n15031), .O(new_n17059));
  nor2 g16866(.a(new_n17059), .b(new_n17056), .O(new_n17060));
  inv1 g16867(.a(new_n17060), .O(new_n17061));
  nor2 g16868(.a(new_n17061), .b(new_n17055), .O(new_n17062));
  inv1 g16869(.a(new_n17055), .O(new_n17063));
  nor2 g16870(.a(new_n17060), .b(new_n17063), .O(new_n17064));
  nor2 g16871(.a(new_n17064), .b(new_n17062), .O(new_n17065));
  nor2 g16872(.a(new_n8946), .b(new_n1903), .O(new_n17066));
  inv1 g16873(.a(new_n17066), .O(new_n17067));
  nor2 g16874(.a(new_n5178), .b(new_n4366), .O(new_n17068));
  nor2 g16875(.a(new_n5393), .b(new_n4093), .O(new_n17069));
  nor2 g16876(.a(new_n17069), .b(new_n17068), .O(new_n17070));
  nor2 g16877(.a(new_n5393), .b(new_n4366), .O(new_n17071));
  inv1 g16878(.a(new_n17071), .O(new_n17072));
  nor2 g16879(.a(new_n17072), .b(new_n16822), .O(new_n17073));
  nor2 g16880(.a(new_n17073), .b(new_n17070), .O(new_n17074));
  nor2 g16881(.a(new_n17074), .b(new_n17067), .O(new_n17075));
  inv1 g16882(.a(new_n17074), .O(new_n17076));
  nor2 g16883(.a(new_n17076), .b(new_n17066), .O(new_n17077));
  nor2 g16884(.a(new_n17077), .b(new_n17075), .O(new_n17078));
  nor2 g16885(.a(new_n17078), .b(new_n17065), .O(new_n17079));
  inv1 g16886(.a(new_n17065), .O(new_n17080));
  inv1 g16887(.a(new_n17078), .O(new_n17081));
  nor2 g16888(.a(new_n17081), .b(new_n17080), .O(new_n17082));
  nor2 g16889(.a(new_n17082), .b(new_n17079), .O(new_n17083));
  nor2 g16890(.a(new_n17083), .b(new_n17054), .O(new_n17084));
  inv1 g16891(.a(new_n17083), .O(new_n17085));
  nor2 g16892(.a(new_n17085), .b(new_n17053), .O(new_n17086));
  nor2 g16893(.a(new_n17086), .b(new_n17084), .O(new_n17087));
  inv1 g16894(.a(new_n17087), .O(new_n17088));
  nor2 g16895(.a(new_n17088), .b(new_n17041), .O(new_n17089));
  nor2 g16896(.a(new_n17087), .b(new_n17040), .O(new_n17090));
  nor2 g16897(.a(new_n17090), .b(new_n17089), .O(new_n17091));
  inv1 g16898(.a(new_n17091), .O(new_n17092));
  nor2 g16899(.a(new_n17092), .b(new_n17005), .O(new_n17093));
  nor2 g16900(.a(new_n17091), .b(new_n17004), .O(new_n17094));
  nor2 g16901(.a(new_n17094), .b(new_n17093), .O(new_n17095));
  inv1 g16902(.a(new_n17095), .O(new_n17096));
  nor2 g16903(.a(new_n17096), .b(new_n16959), .O(new_n17097));
  inv1 g16904(.a(new_n16959), .O(new_n17098));
  nor2 g16905(.a(new_n17095), .b(new_n17098), .O(new_n17099));
  nor2 g16906(.a(new_n17099), .b(new_n17097), .O(new_n17100));
  inv1 g16907(.a(new_n17100), .O(new_n17101));
  nor2 g16908(.a(new_n17101), .b(new_n16958), .O(new_n17102));
  inv1 g16909(.a(new_n16958), .O(new_n17103));
  nor2 g16910(.a(new_n17100), .b(new_n17103), .O(new_n17104));
  nor2 g16911(.a(new_n17104), .b(new_n17102), .O(new_n17105));
  nor2 g16912(.a(new_n17105), .b(new_n16957), .O(new_n17106));
  inv1 g16913(.a(new_n17105), .O(new_n17107));
  nor2 g16914(.a(new_n17107), .b(new_n16956), .O(new_n17108));
  nor2 g16915(.a(new_n17108), .b(new_n17106), .O(new_n17109));
  inv1 g16916(.a(new_n17109), .O(new_n17110));
  nor2 g16917(.a(new_n16929), .b(new_n16900), .O(new_n17111));
  nor2 g16918(.a(new_n16894), .b(new_n16891), .O(new_n17112));
  nor2 g16919(.a(new_n16706), .b(new_n16699), .O(new_n17113));
  nor2 g16920(.a(new_n16817), .b(new_n16811), .O(new_n17114));
  nor2 g16921(.a(new_n17114), .b(new_n17113), .O(new_n17115));
  inv1 g16922(.a(new_n17113), .O(new_n17116));
  inv1 g16923(.a(new_n17114), .O(new_n17117));
  nor2 g16924(.a(new_n17117), .b(new_n17116), .O(new_n17118));
  nor2 g16925(.a(new_n17118), .b(new_n17115), .O(new_n17119));
  nor2 g16926(.a(new_n16719), .b(new_n16712), .O(new_n17120));
  nor2 g16927(.a(new_n17120), .b(new_n17119), .O(new_n17121));
  inv1 g16928(.a(new_n17119), .O(new_n17122));
  inv1 g16929(.a(new_n17120), .O(new_n17123));
  nor2 g16930(.a(new_n17123), .b(new_n17122), .O(new_n17124));
  nor2 g16931(.a(new_n17124), .b(new_n17121), .O(new_n17125));
  nor2 g16932(.a(new_n16728), .b(new_n16721), .O(new_n17126));
  inv1 g16933(.a(new_n17126), .O(new_n17127));
  nor2 g16934(.a(new_n17127), .b(new_n17125), .O(new_n17128));
  inv1 g16935(.a(new_n17125), .O(new_n17129));
  nor2 g16936(.a(new_n17126), .b(new_n17129), .O(new_n17130));
  nor2 g16937(.a(new_n17130), .b(new_n17128), .O(new_n17131));
  nor2 g16938(.a(new_n16914), .b(new_n16908), .O(new_n17132));
  inv1 g16939(.a(new_n17132), .O(new_n17133));
  nor2 g16940(.a(new_n17133), .b(new_n17131), .O(new_n17134));
  inv1 g16941(.a(new_n17131), .O(new_n17135));
  nor2 g16942(.a(new_n17132), .b(new_n17135), .O(new_n17136));
  nor2 g16943(.a(new_n17136), .b(new_n17134), .O(new_n17137));
  inv1 g16944(.a(new_n17137), .O(new_n17138));
  nor2 g16945(.a(new_n17138), .b(new_n17112), .O(new_n17139));
  inv1 g16946(.a(new_n17112), .O(new_n17140));
  nor2 g16947(.a(new_n17137), .b(new_n17140), .O(new_n17141));
  nor2 g16948(.a(new_n17141), .b(new_n17139), .O(new_n17142));
  inv1 g16949(.a(new_n17142), .O(new_n17143));
  nor2 g16950(.a(new_n16877), .b(new_n16870), .O(new_n17144));
  nor2 g16951(.a(new_n16863), .b(new_n16859), .O(new_n17145));
  nor2 g16952(.a(new_n17145), .b(new_n17144), .O(new_n17146));
  inv1 g16953(.a(new_n17144), .O(new_n17147));
  inv1 g16954(.a(new_n17145), .O(new_n17148));
  nor2 g16955(.a(new_n17148), .b(new_n17147), .O(new_n17149));
  nor2 g16956(.a(new_n17149), .b(new_n17146), .O(new_n17150));
  nor2 g16957(.a(new_n16853), .b(new_n16846), .O(new_n17151));
  nor2 g16958(.a(new_n17151), .b(new_n17150), .O(new_n17152));
  inv1 g16959(.a(new_n17150), .O(new_n17153));
  inv1 g16960(.a(new_n17151), .O(new_n17154));
  nor2 g16961(.a(new_n17154), .b(new_n17153), .O(new_n17155));
  nor2 g16962(.a(new_n17155), .b(new_n17152), .O(new_n17156));
  inv1 g16963(.a(new_n17156), .O(new_n17157));
  nor2 g16964(.a(new_n16840), .b(new_n16834), .O(new_n17158));
  inv1 g16965(.a(new_n17158), .O(new_n17159));
  nor2 g16966(.a(new_n16886), .b(new_n16879), .O(new_n17160));
  inv1 g16967(.a(new_n17160), .O(new_n17161));
  nor2 g16968(.a(new_n17161), .b(new_n17159), .O(new_n17162));
  nor2 g16969(.a(new_n17160), .b(new_n17158), .O(new_n17163));
  nor2 g16970(.a(new_n17163), .b(new_n17162), .O(new_n17164));
  inv1 g16971(.a(new_n17164), .O(new_n17165));
  nor2 g16972(.a(new_n17165), .b(new_n17157), .O(new_n17166));
  nor2 g16973(.a(new_n17164), .b(new_n17156), .O(new_n17167));
  nor2 g16974(.a(new_n17167), .b(new_n17166), .O(new_n17168));
  inv1 g16975(.a(new_n17168), .O(new_n17169));
  nor2 g16976(.a(new_n17169), .b(new_n17143), .O(new_n17170));
  nor2 g16977(.a(new_n17168), .b(new_n17142), .O(new_n17171));
  nor2 g16978(.a(new_n17171), .b(new_n17170), .O(new_n17172));
  inv1 g16979(.a(new_n17172), .O(new_n17173));
  nor2 g16980(.a(new_n16686), .b(new_n16680), .O(new_n17174));
  inv1 g16981(.a(new_n17174), .O(new_n17175));
  nor2 g16982(.a(new_n16764), .b(new_n16758), .O(new_n17176));
  inv1 g16983(.a(new_n17176), .O(new_n17177));
  nor2 g16984(.a(new_n17177), .b(new_n17175), .O(new_n17178));
  nor2 g16985(.a(new_n17176), .b(new_n17174), .O(new_n17179));
  nor2 g16986(.a(new_n17179), .b(new_n17178), .O(new_n17180));
  nor2 g16987(.a(new_n16750), .b(new_n16743), .O(new_n17181));
  inv1 g16988(.a(new_n17181), .O(new_n17182));
  nor2 g16989(.a(new_n17182), .b(new_n17180), .O(new_n17183));
  inv1 g16990(.a(new_n17180), .O(new_n17184));
  nor2 g16991(.a(new_n17181), .b(new_n17184), .O(new_n17185));
  nor2 g16992(.a(new_n17185), .b(new_n17183), .O(new_n17186));
  nor2 g16993(.a(new_n16731), .b(new_n16692), .O(new_n17187));
  nor2 g16994(.a(new_n16772), .b(new_n16767), .O(new_n17188));
  nor2 g16995(.a(new_n17188), .b(new_n17187), .O(new_n17189));
  inv1 g16996(.a(new_n17187), .O(new_n17190));
  inv1 g16997(.a(new_n17188), .O(new_n17191));
  nor2 g16998(.a(new_n17191), .b(new_n17190), .O(new_n17192));
  nor2 g16999(.a(new_n17192), .b(new_n17189), .O(new_n17193));
  nor2 g17000(.a(new_n17193), .b(new_n17186), .O(new_n17194));
  inv1 g17001(.a(new_n17186), .O(new_n17195));
  inv1 g17002(.a(new_n17193), .O(new_n17196));
  nor2 g17003(.a(new_n17196), .b(new_n17195), .O(new_n17197));
  nor2 g17004(.a(new_n17197), .b(new_n17194), .O(new_n17198));
  inv1 g17005(.a(new_n17198), .O(new_n17199));
  nor2 g17006(.a(new_n17199), .b(new_n17173), .O(new_n17200));
  nor2 g17007(.a(new_n17198), .b(new_n17172), .O(new_n17201));
  nor2 g17008(.a(new_n17201), .b(new_n17200), .O(new_n17202));
  inv1 g17009(.a(new_n17202), .O(new_n17203));
  nor2 g17010(.a(new_n17203), .b(new_n17111), .O(new_n17204));
  inv1 g17011(.a(new_n17111), .O(new_n17205));
  nor2 g17012(.a(new_n17202), .b(new_n17205), .O(new_n17206));
  nor2 g17013(.a(new_n17206), .b(new_n17204), .O(new_n17207));
  inv1 g17014(.a(new_n17207), .O(new_n17208));
  nor2 g17015(.a(new_n17208), .b(new_n17110), .O(new_n17209));
  nor2 g17016(.a(new_n17207), .b(new_n17109), .O(new_n17210));
  nor2 g17017(.a(new_n17210), .b(new_n17209), .O(new_n17211));
  nor2 g17018(.a(new_n17211), .b(new_n16955), .O(new_n17212));
  inv1 g17019(.a(new_n17211), .O(new_n17213));
  nor2 g17020(.a(new_n17213), .b(new_n16954), .O(new_n17214));
  nor2 g17021(.a(new_n17214), .b(new_n17212), .O(new_n17215));
  inv1 g17022(.a(new_n17215), .O(new_n17216));
  nor2 g17023(.a(new_n16949), .b(new_n16945), .O(new_n17217));
  nor2 g17024(.a(new_n17217), .b(new_n17216), .O(new_n17218));
  inv1 g17025(.a(new_n17217), .O(new_n17219));
  nor2 g17026(.a(new_n17219), .b(new_n17215), .O(new_n17220));
  nor2 g17027(.a(new_n17220), .b(new_n17218), .O(new_n17221));
  inv1 g17028(.a(new_n17221), .O(\asquared[81] ));
  nor2 g17029(.a(new_n17209), .b(new_n17108), .O(new_n17223));
  nor2 g17030(.a(new_n17204), .b(new_n17200), .O(new_n17224));
  nor2 g17031(.a(new_n17170), .b(new_n17139), .O(new_n17225));
  nor2 g17032(.a(new_n17197), .b(new_n17189), .O(new_n17226));
  nor2 g17033(.a(new_n17185), .b(new_n17179), .O(new_n17227));
  inv1 g17034(.a(new_n17227), .O(new_n17228));
  nor2 g17035(.a(new_n6893), .b(new_n3231), .O(new_n17229));
  nor2 g17036(.a(new_n6570), .b(new_n3533), .O(new_n17230));
  nor2 g17037(.a(new_n17230), .b(new_n17229), .O(new_n17231));
  nor2 g17038(.a(new_n6893), .b(new_n3533), .O(new_n17232));
  inv1 g17039(.a(new_n17232), .O(new_n17233));
  nor2 g17040(.a(new_n17233), .b(new_n16848), .O(new_n17234));
  nor2 g17041(.a(new_n17234), .b(new_n17231), .O(new_n17235));
  nor2 g17042(.a(new_n17235), .b(new_n12580), .O(new_n17236));
  inv1 g17043(.a(new_n17235), .O(new_n17237));
  nor2 g17044(.a(new_n17237), .b(new_n12579), .O(new_n17238));
  nor2 g17045(.a(new_n17238), .b(new_n17236), .O(new_n17239));
  inv1 g17046(.a(new_n17239), .O(new_n17240));
  nor2 g17047(.a(new_n9873), .b(new_n1647), .O(new_n17241));
  nor2 g17048(.a(new_n17241), .b(new_n15409), .O(new_n17242));
  inv1 g17049(.a(new_n16710), .O(new_n17243));
  nor2 g17050(.a(new_n9873), .b(new_n1903), .O(new_n17244));
  inv1 g17051(.a(new_n17244), .O(new_n17245));
  nor2 g17052(.a(new_n17245), .b(new_n17243), .O(new_n17246));
  nor2 g17053(.a(new_n17246), .b(new_n17242), .O(new_n17247));
  nor2 g17054(.a(new_n17247), .b(new_n17010), .O(new_n17248));
  inv1 g17055(.a(new_n17247), .O(new_n17249));
  nor2 g17056(.a(new_n17249), .b(new_n17009), .O(new_n17250));
  nor2 g17057(.a(new_n17250), .b(new_n17248), .O(new_n17251));
  nor2 g17058(.a(new_n4954), .b(\a[40] ), .O(new_n17252));
  nor2 g17059(.a(new_n17252), .b(new_n16964), .O(new_n17253));
  inv1 g17060(.a(new_n17252), .O(new_n17254));
  nor2 g17061(.a(new_n17254), .b(new_n16963), .O(new_n17255));
  nor2 g17062(.a(new_n17255), .b(new_n17253), .O(new_n17256));
  nor2 g17063(.a(new_n17256), .b(new_n17251), .O(new_n17257));
  inv1 g17064(.a(new_n17251), .O(new_n17258));
  inv1 g17065(.a(new_n17256), .O(new_n17259));
  nor2 g17066(.a(new_n17259), .b(new_n17258), .O(new_n17260));
  nor2 g17067(.a(new_n17260), .b(new_n17257), .O(new_n17261));
  nor2 g17068(.a(new_n17261), .b(new_n17240), .O(new_n17262));
  inv1 g17069(.a(new_n17261), .O(new_n17263));
  nor2 g17070(.a(new_n17263), .b(new_n17239), .O(new_n17264));
  nor2 g17071(.a(new_n17264), .b(new_n17262), .O(new_n17265));
  nor2 g17072(.a(new_n17265), .b(new_n17228), .O(new_n17266));
  inv1 g17073(.a(new_n17265), .O(new_n17267));
  nor2 g17074(.a(new_n17267), .b(new_n17227), .O(new_n17268));
  nor2 g17075(.a(new_n17268), .b(new_n17266), .O(new_n17269));
  nor2 g17076(.a(new_n11596), .b(new_n1086), .O(new_n17270));
  nor2 g17077(.a(new_n10895), .b(new_n1297), .O(new_n17271));
  nor2 g17078(.a(new_n10468), .b(new_n1425), .O(new_n17272));
  nor2 g17079(.a(new_n17272), .b(new_n17271), .O(new_n17273));
  nor2 g17080(.a(new_n10895), .b(new_n1425), .O(new_n17274));
  inv1 g17081(.a(new_n17274), .O(new_n17275));
  nor2 g17082(.a(new_n17275), .b(new_n17016), .O(new_n17276));
  nor2 g17083(.a(new_n17276), .b(new_n17273), .O(new_n17277));
  inv1 g17084(.a(new_n17277), .O(new_n17278));
  nor2 g17085(.a(new_n17278), .b(new_n17270), .O(new_n17279));
  inv1 g17086(.a(new_n17270), .O(new_n17280));
  nor2 g17087(.a(new_n17277), .b(new_n17280), .O(new_n17281));
  nor2 g17088(.a(new_n17281), .b(new_n17279), .O(new_n17282));
  nor2 g17089(.a(new_n6274), .b(new_n3722), .O(new_n17283));
  inv1 g17090(.a(new_n17283), .O(new_n17284));
  nor2 g17091(.a(new_n5796), .b(new_n4093), .O(new_n17285));
  nor2 g17092(.a(new_n17285), .b(new_n16988), .O(new_n17286));
  inv1 g17093(.a(new_n16985), .O(new_n17287));
  nor2 g17094(.a(new_n5971), .b(new_n4093), .O(new_n17288));
  inv1 g17095(.a(new_n17288), .O(new_n17289));
  nor2 g17096(.a(new_n17289), .b(new_n17287), .O(new_n17290));
  nor2 g17097(.a(new_n17290), .b(new_n17286), .O(new_n17291));
  nor2 g17098(.a(new_n17291), .b(new_n17284), .O(new_n17292));
  inv1 g17099(.a(new_n17291), .O(new_n17293));
  nor2 g17100(.a(new_n17293), .b(new_n17283), .O(new_n17294));
  nor2 g17101(.a(new_n17294), .b(new_n17292), .O(new_n17295));
  nor2 g17102(.a(new_n17295), .b(new_n17282), .O(new_n17296));
  inv1 g17103(.a(new_n17282), .O(new_n17297));
  inv1 g17104(.a(new_n17295), .O(new_n17298));
  nor2 g17105(.a(new_n17298), .b(new_n17297), .O(new_n17299));
  nor2 g17106(.a(new_n17299), .b(new_n17296), .O(new_n17300));
  inv1 g17107(.a(new_n17300), .O(new_n17301));
  nor2 g17108(.a(new_n8946), .b(new_n2121), .O(new_n17302));
  inv1 g17109(.a(new_n17302), .O(new_n17303));
  nor2 g17110(.a(new_n8026), .b(new_n2506), .O(new_n17304));
  nor2 g17111(.a(new_n17304), .b(new_n17046), .O(new_n17305));
  inv1 g17112(.a(new_n17043), .O(new_n17306));
  nor2 g17113(.a(new_n8170), .b(new_n2506), .O(new_n17307));
  inv1 g17114(.a(new_n17307), .O(new_n17308));
  nor2 g17115(.a(new_n17308), .b(new_n17306), .O(new_n17309));
  nor2 g17116(.a(new_n17309), .b(new_n17305), .O(new_n17310));
  nor2 g17117(.a(new_n17310), .b(new_n17303), .O(new_n17311));
  inv1 g17118(.a(new_n17310), .O(new_n17312));
  nor2 g17119(.a(new_n17312), .b(new_n17302), .O(new_n17313));
  nor2 g17120(.a(new_n17313), .b(new_n17311), .O(new_n17314));
  nor2 g17121(.a(new_n17314), .b(new_n17301), .O(new_n17315));
  inv1 g17122(.a(new_n17314), .O(new_n17316));
  nor2 g17123(.a(new_n17316), .b(new_n17300), .O(new_n17317));
  nor2 g17124(.a(new_n17317), .b(new_n17315), .O(new_n17318));
  nor2 g17125(.a(new_n17318), .b(new_n17269), .O(new_n17319));
  inv1 g17126(.a(new_n17269), .O(new_n17320));
  inv1 g17127(.a(new_n17318), .O(new_n17321));
  nor2 g17128(.a(new_n17321), .b(new_n17320), .O(new_n17322));
  nor2 g17129(.a(new_n17322), .b(new_n17319), .O(new_n17323));
  inv1 g17130(.a(new_n17323), .O(new_n17324));
  nor2 g17131(.a(new_n17324), .b(new_n17226), .O(new_n17325));
  inv1 g17132(.a(new_n17226), .O(new_n17326));
  nor2 g17133(.a(new_n17323), .b(new_n17326), .O(new_n17327));
  nor2 g17134(.a(new_n17327), .b(new_n17325), .O(new_n17328));
  inv1 g17135(.a(new_n17328), .O(new_n17329));
  nor2 g17136(.a(new_n17329), .b(new_n17225), .O(new_n17330));
  inv1 g17137(.a(new_n17225), .O(new_n17331));
  nor2 g17138(.a(new_n17328), .b(new_n17331), .O(new_n17332));
  nor2 g17139(.a(new_n17332), .b(new_n17330), .O(new_n17333));
  inv1 g17140(.a(new_n17333), .O(new_n17334));
  nor2 g17141(.a(new_n17334), .b(new_n17224), .O(new_n17335));
  inv1 g17142(.a(new_n17224), .O(new_n17336));
  nor2 g17143(.a(new_n17333), .b(new_n17336), .O(new_n17337));
  nor2 g17144(.a(new_n17337), .b(new_n17335), .O(new_n17338));
  inv1 g17145(.a(new_n17338), .O(new_n17339));
  nor2 g17146(.a(new_n17093), .b(new_n17089), .O(new_n17340));
  inv1 g17147(.a(new_n17340), .O(new_n17341));
  nor2 g17148(.a(new_n17035), .b(new_n17028), .O(new_n17342));
  nor2 g17149(.a(new_n16980), .b(new_n16974), .O(new_n17343));
  nor2 g17150(.a(new_n17343), .b(new_n17342), .O(new_n17344));
  inv1 g17151(.a(new_n17342), .O(new_n17345));
  inv1 g17152(.a(new_n17343), .O(new_n17346));
  nor2 g17153(.a(new_n17346), .b(new_n17345), .O(new_n17347));
  nor2 g17154(.a(new_n17347), .b(new_n17344), .O(new_n17348));
  nor2 g17155(.a(new_n17017), .b(new_n17011), .O(new_n17349));
  inv1 g17156(.a(new_n17349), .O(new_n17350));
  nor2 g17157(.a(new_n17350), .b(new_n17348), .O(new_n17351));
  inv1 g17158(.a(new_n17348), .O(new_n17352));
  nor2 g17159(.a(new_n17349), .b(new_n17352), .O(new_n17353));
  nor2 g17160(.a(new_n17353), .b(new_n17351), .O(new_n17354));
  inv1 g17161(.a(new_n17354), .O(new_n17355));
  nor2 g17162(.a(new_n17002), .b(new_n16996), .O(new_n17356));
  nor2 g17163(.a(new_n17356), .b(new_n17355), .O(new_n17357));
  inv1 g17164(.a(new_n17356), .O(new_n17358));
  nor2 g17165(.a(new_n17358), .b(new_n17354), .O(new_n17359));
  nor2 g17166(.a(new_n17359), .b(new_n17357), .O(new_n17360));
  inv1 g17167(.a(new_n17360), .O(new_n17361));
  nor2 g17168(.a(new_n16968), .b(new_n16965), .O(new_n17362));
  inv1 g17169(.a(new_n17362), .O(new_n17363));
  nor2 g17170(.a(new_n16994), .b(new_n16986), .O(new_n17364));
  nor2 g17171(.a(new_n17364), .b(new_n17363), .O(new_n17365));
  inv1 g17172(.a(new_n17364), .O(new_n17366));
  nor2 g17173(.a(new_n17366), .b(new_n17362), .O(new_n17367));
  nor2 g17174(.a(new_n17367), .b(new_n17365), .O(new_n17368));
  inv1 g17175(.a(new_n17368), .O(new_n17369));
  nor2 g17176(.a(new_n7537), .b(new_n2660), .O(new_n17370));
  inv1 g17177(.a(new_n17370), .O(new_n17371));
  nor2 g17178(.a(new_n7294), .b(new_n2826), .O(new_n17372));
  nor2 g17179(.a(new_n17372), .b(new_n17029), .O(new_n17373));
  inv1 g17180(.a(new_n17026), .O(new_n17374));
  nor2 g17181(.a(new_n7294), .b(new_n3057), .O(new_n17375));
  inv1 g17182(.a(new_n17375), .O(new_n17376));
  nor2 g17183(.a(new_n17376), .b(new_n17374), .O(new_n17377));
  nor2 g17184(.a(new_n17377), .b(new_n17373), .O(new_n17378));
  nor2 g17185(.a(new_n17378), .b(new_n17371), .O(new_n17379));
  inv1 g17186(.a(new_n17378), .O(new_n17380));
  nor2 g17187(.a(new_n17380), .b(new_n17370), .O(new_n17381));
  nor2 g17188(.a(new_n17381), .b(new_n17379), .O(new_n17382));
  nor2 g17189(.a(new_n17382), .b(new_n17369), .O(new_n17383));
  inv1 g17190(.a(new_n17382), .O(new_n17384));
  nor2 g17191(.a(new_n17384), .b(new_n17368), .O(new_n17385));
  nor2 g17192(.a(new_n17385), .b(new_n17383), .O(new_n17386));
  inv1 g17193(.a(new_n17386), .O(new_n17387));
  nor2 g17194(.a(new_n17387), .b(new_n17361), .O(new_n17388));
  nor2 g17195(.a(new_n17386), .b(new_n17360), .O(new_n17389));
  nor2 g17196(.a(new_n17389), .b(new_n17388), .O(new_n17390));
  nor2 g17197(.a(new_n17390), .b(new_n17341), .O(new_n17391));
  inv1 g17198(.a(new_n17390), .O(new_n17392));
  nor2 g17199(.a(new_n17392), .b(new_n17340), .O(new_n17393));
  nor2 g17200(.a(new_n17393), .b(new_n17391), .O(new_n17394));
  inv1 g17201(.a(new_n17394), .O(new_n17395));
  nor2 g17202(.a(new_n17077), .b(new_n17070), .O(new_n17396));
  nor2 g17203(.a(new_n17052), .b(new_n17044), .O(new_n17397));
  nor2 g17204(.a(new_n17397), .b(new_n17396), .O(new_n17398));
  inv1 g17205(.a(new_n17396), .O(new_n17399));
  inv1 g17206(.a(new_n17397), .O(new_n17400));
  nor2 g17207(.a(new_n17400), .b(new_n17399), .O(new_n17401));
  nor2 g17208(.a(new_n17401), .b(new_n17398), .O(new_n17402));
  nor2 g17209(.a(new_n17062), .b(new_n17056), .O(new_n17403));
  nor2 g17210(.a(new_n17403), .b(new_n17402), .O(new_n17404));
  inv1 g17211(.a(new_n17402), .O(new_n17405));
  inv1 g17212(.a(new_n17403), .O(new_n17406));
  nor2 g17213(.a(new_n17406), .b(new_n17405), .O(new_n17407));
  nor2 g17214(.a(new_n17407), .b(new_n17404), .O(new_n17408));
  inv1 g17215(.a(new_n17408), .O(new_n17409));
  nor2 g17216(.a(new_n17037), .b(new_n17022), .O(new_n17410));
  inv1 g17217(.a(new_n17410), .O(new_n17411));
  nor2 g17218(.a(new_n17086), .b(new_n17079), .O(new_n17412));
  inv1 g17219(.a(new_n17412), .O(new_n17413));
  nor2 g17220(.a(new_n17413), .b(new_n17411), .O(new_n17414));
  nor2 g17221(.a(new_n17412), .b(new_n17410), .O(new_n17415));
  nor2 g17222(.a(new_n17415), .b(new_n17414), .O(new_n17416));
  inv1 g17223(.a(new_n17416), .O(new_n17417));
  nor2 g17224(.a(new_n17417), .b(new_n17409), .O(new_n17418));
  nor2 g17225(.a(new_n17416), .b(new_n17408), .O(new_n17419));
  nor2 g17226(.a(new_n17419), .b(new_n17418), .O(new_n17420));
  inv1 g17227(.a(new_n17420), .O(new_n17421));
  nor2 g17228(.a(new_n17421), .b(new_n17395), .O(new_n17422));
  nor2 g17229(.a(new_n17420), .b(new_n17394), .O(new_n17423));
  nor2 g17230(.a(new_n17423), .b(new_n17422), .O(new_n17424));
  inv1 g17231(.a(new_n17424), .O(new_n17425));
  nor2 g17232(.a(new_n17102), .b(new_n17097), .O(new_n17426));
  nor2 g17233(.a(new_n17124), .b(new_n17118), .O(new_n17427));
  inv1 g17234(.a(new_n17427), .O(new_n17428));
  nor2 g17235(.a(new_n17155), .b(new_n17149), .O(new_n17429));
  nor2 g17236(.a(new_n8476), .b(new_n2184), .O(new_n17430));
  inv1 g17237(.a(new_n17430), .O(new_n17431));
  nor2 g17238(.a(new_n5178), .b(new_n4425), .O(new_n17432));
  nor2 g17239(.a(new_n17432), .b(new_n17071), .O(new_n17433));
  inv1 g17240(.a(new_n17068), .O(new_n17434));
  nor2 g17241(.a(new_n5393), .b(new_n4425), .O(new_n17435));
  inv1 g17242(.a(new_n17435), .O(new_n17436));
  nor2 g17243(.a(new_n17436), .b(new_n17434), .O(new_n17437));
  nor2 g17244(.a(new_n17437), .b(new_n17433), .O(new_n17438));
  nor2 g17245(.a(new_n17438), .b(new_n17431), .O(new_n17439));
  inv1 g17246(.a(new_n17438), .O(new_n17440));
  nor2 g17247(.a(new_n17440), .b(new_n17430), .O(new_n17441));
  nor2 g17248(.a(new_n17441), .b(new_n17439), .O(new_n17442));
  nor2 g17249(.a(new_n17442), .b(new_n17429), .O(new_n17443));
  inv1 g17250(.a(new_n17429), .O(new_n17444));
  inv1 g17251(.a(new_n17442), .O(new_n17445));
  nor2 g17252(.a(new_n17445), .b(new_n17444), .O(new_n17446));
  nor2 g17253(.a(new_n17446), .b(new_n17443), .O(new_n17447));
  nor2 g17254(.a(new_n17447), .b(new_n17428), .O(new_n17448));
  inv1 g17255(.a(new_n17447), .O(new_n17449));
  nor2 g17256(.a(new_n17449), .b(new_n17427), .O(new_n17450));
  nor2 g17257(.a(new_n17450), .b(new_n17448), .O(new_n17451));
  inv1 g17258(.a(new_n17451), .O(new_n17452));
  nor2 g17259(.a(new_n17136), .b(new_n17130), .O(new_n17453));
  nor2 g17260(.a(new_n17166), .b(new_n17163), .O(new_n17454));
  nor2 g17261(.a(new_n17454), .b(new_n17453), .O(new_n17455));
  inv1 g17262(.a(new_n17453), .O(new_n17456));
  inv1 g17263(.a(new_n17454), .O(new_n17457));
  nor2 g17264(.a(new_n17457), .b(new_n17456), .O(new_n17458));
  nor2 g17265(.a(new_n17458), .b(new_n17455), .O(new_n17459));
  inv1 g17266(.a(new_n17459), .O(new_n17460));
  nor2 g17267(.a(new_n17460), .b(new_n17452), .O(new_n17461));
  nor2 g17268(.a(new_n17459), .b(new_n17451), .O(new_n17462));
  nor2 g17269(.a(new_n17462), .b(new_n17461), .O(new_n17463));
  inv1 g17270(.a(new_n17463), .O(new_n17464));
  nor2 g17271(.a(new_n17464), .b(new_n17426), .O(new_n17465));
  inv1 g17272(.a(new_n17426), .O(new_n17466));
  nor2 g17273(.a(new_n17463), .b(new_n17466), .O(new_n17467));
  nor2 g17274(.a(new_n17467), .b(new_n17465), .O(new_n17468));
  inv1 g17275(.a(new_n17468), .O(new_n17469));
  nor2 g17276(.a(new_n17469), .b(new_n17425), .O(new_n17470));
  nor2 g17277(.a(new_n17468), .b(new_n17424), .O(new_n17471));
  nor2 g17278(.a(new_n17471), .b(new_n17470), .O(new_n17472));
  inv1 g17279(.a(new_n17472), .O(new_n17473));
  nor2 g17280(.a(new_n17473), .b(new_n17339), .O(new_n17474));
  nor2 g17281(.a(new_n17472), .b(new_n17338), .O(new_n17475));
  nor2 g17282(.a(new_n17475), .b(new_n17474), .O(new_n17476));
  inv1 g17283(.a(new_n17476), .O(new_n17477));
  nor2 g17284(.a(new_n17477), .b(new_n17223), .O(new_n17478));
  inv1 g17285(.a(new_n17223), .O(new_n17479));
  nor2 g17286(.a(new_n17476), .b(new_n17479), .O(new_n17480));
  nor2 g17287(.a(new_n17480), .b(new_n17478), .O(new_n17481));
  inv1 g17288(.a(new_n17481), .O(new_n17482));
  nor2 g17289(.a(new_n17218), .b(new_n17212), .O(new_n17483));
  nor2 g17290(.a(new_n17483), .b(new_n17482), .O(new_n17484));
  inv1 g17291(.a(new_n17483), .O(new_n17485));
  nor2 g17292(.a(new_n17485), .b(new_n17481), .O(new_n17486));
  nor2 g17293(.a(new_n17486), .b(new_n17484), .O(new_n17487));
  inv1 g17294(.a(new_n17487), .O(\asquared[82] ));
  nor2 g17295(.a(new_n17474), .b(new_n17335), .O(new_n17489));
  nor2 g17296(.a(new_n17470), .b(new_n17465), .O(new_n17490));
  nor2 g17297(.a(new_n17422), .b(new_n17393), .O(new_n17491));
  nor2 g17298(.a(new_n17461), .b(new_n17455), .O(new_n17492));
  nor2 g17299(.a(new_n17450), .b(new_n17443), .O(new_n17493));
  inv1 g17300(.a(new_n17493), .O(new_n17494));
  nor2 g17301(.a(new_n10468), .b(new_n1493), .O(new_n17495));
  inv1 g17302(.a(new_n17495), .O(new_n17496));
  nor2 g17303(.a(new_n9873), .b(new_n1736), .O(new_n17497));
  nor2 g17304(.a(new_n10320), .b(new_n1647), .O(new_n17498));
  nor2 g17305(.a(new_n17498), .b(new_n17497), .O(new_n17499));
  inv1 g17306(.a(new_n17241), .O(new_n17500));
  nor2 g17307(.a(new_n10320), .b(new_n1736), .O(new_n17501));
  inv1 g17308(.a(new_n17501), .O(new_n17502));
  nor2 g17309(.a(new_n17502), .b(new_n17500), .O(new_n17503));
  nor2 g17310(.a(new_n17503), .b(new_n17499), .O(new_n17504));
  nor2 g17311(.a(new_n17504), .b(new_n17496), .O(new_n17505));
  inv1 g17312(.a(new_n17504), .O(new_n17506));
  nor2 g17313(.a(new_n17506), .b(new_n17495), .O(new_n17507));
  nor2 g17314(.a(new_n17507), .b(new_n17505), .O(new_n17508));
  inv1 g17315(.a(new_n17508), .O(new_n17509));
  nor2 g17316(.a(new_n6958), .b(new_n3231), .O(new_n17510));
  nor2 g17317(.a(new_n17510), .b(new_n17232), .O(new_n17511));
  inv1 g17318(.a(new_n17229), .O(new_n17512));
  nor2 g17319(.a(new_n6958), .b(new_n3533), .O(new_n17513));
  inv1 g17320(.a(new_n17513), .O(new_n17514));
  nor2 g17321(.a(new_n17514), .b(new_n17512), .O(new_n17515));
  nor2 g17322(.a(new_n17515), .b(new_n17511), .O(new_n17516));
  nor2 g17323(.a(new_n17516), .b(new_n17376), .O(new_n17517));
  inv1 g17324(.a(new_n17516), .O(new_n17518));
  nor2 g17325(.a(new_n17518), .b(new_n17375), .O(new_n17519));
  nor2 g17326(.a(new_n17519), .b(new_n17517), .O(new_n17520));
  nor2 g17327(.a(new_n11186), .b(new_n1297), .O(new_n17521));
  inv1 g17328(.a(new_n17521), .O(new_n17522));
  nor2 g17329(.a(new_n7537), .b(new_n2826), .O(new_n17523));
  nor2 g17330(.a(new_n17523), .b(new_n17274), .O(new_n17524));
  inv1 g17331(.a(new_n17523), .O(new_n17525));
  nor2 g17332(.a(new_n17525), .b(new_n17275), .O(new_n17526));
  nor2 g17333(.a(new_n17526), .b(new_n17524), .O(new_n17527));
  nor2 g17334(.a(new_n17527), .b(new_n17522), .O(new_n17528));
  inv1 g17335(.a(new_n17527), .O(new_n17529));
  nor2 g17336(.a(new_n17529), .b(new_n17521), .O(new_n17530));
  nor2 g17337(.a(new_n17530), .b(new_n17528), .O(new_n17531));
  nor2 g17338(.a(new_n17531), .b(new_n17520), .O(new_n17532));
  inv1 g17339(.a(new_n17520), .O(new_n17533));
  inv1 g17340(.a(new_n17531), .O(new_n17534));
  nor2 g17341(.a(new_n17534), .b(new_n17533), .O(new_n17535));
  nor2 g17342(.a(new_n17535), .b(new_n17532), .O(new_n17536));
  nor2 g17343(.a(new_n17536), .b(new_n17509), .O(new_n17537));
  inv1 g17344(.a(new_n17536), .O(new_n17538));
  nor2 g17345(.a(new_n17538), .b(new_n17508), .O(new_n17539));
  nor2 g17346(.a(new_n17539), .b(new_n17537), .O(new_n17540));
  nor2 g17347(.a(new_n17540), .b(new_n17494), .O(new_n17541));
  inv1 g17348(.a(new_n17540), .O(new_n17542));
  nor2 g17349(.a(new_n17542), .b(new_n17493), .O(new_n17543));
  nor2 g17350(.a(new_n17543), .b(new_n17541), .O(new_n17544));
  nor2 g17351(.a(new_n6570), .b(new_n3722), .O(new_n17545));
  inv1 g17352(.a(new_n17545), .O(new_n17546));
  nor2 g17353(.a(new_n6274), .b(new_n3870), .O(new_n17547));
  nor2 g17354(.a(new_n17547), .b(new_n17288), .O(new_n17548));
  nor2 g17355(.a(new_n6274), .b(new_n4093), .O(new_n17549));
  inv1 g17356(.a(new_n17549), .O(new_n17550));
  nor2 g17357(.a(new_n17550), .b(new_n16989), .O(new_n17551));
  nor2 g17358(.a(new_n17551), .b(new_n17548), .O(new_n17552));
  nor2 g17359(.a(new_n17552), .b(new_n17546), .O(new_n17553));
  inv1 g17360(.a(new_n17552), .O(new_n17554));
  nor2 g17361(.a(new_n17554), .b(new_n17545), .O(new_n17555));
  nor2 g17362(.a(new_n17555), .b(new_n17553), .O(new_n17556));
  inv1 g17363(.a(new_n17556), .O(new_n17557));
  nor2 g17364(.a(new_n5796), .b(new_n4366), .O(new_n17558));
  nor2 g17365(.a(new_n17558), .b(new_n17435), .O(new_n17559));
  nor2 g17366(.a(new_n5796), .b(new_n4425), .O(new_n17560));
  inv1 g17367(.a(new_n17560), .O(new_n17561));
  nor2 g17368(.a(new_n17561), .b(new_n17072), .O(new_n17562));
  nor2 g17369(.a(new_n17562), .b(new_n17559), .O(new_n17563));
  inv1 g17370(.a(new_n17563), .O(new_n17564));
  nor2 g17371(.a(new_n17564), .b(new_n17057), .O(new_n17565));
  nor2 g17372(.a(new_n17563), .b(new_n17058), .O(new_n17566));
  nor2 g17373(.a(new_n17566), .b(new_n17565), .O(new_n17567));
  nor2 g17374(.a(new_n5178), .b(new_n4682), .O(new_n17568));
  inv1 g17375(.a(new_n17568), .O(new_n17569));
  nor2 g17376(.a(new_n8026), .b(new_n2660), .O(new_n17570));
  nor2 g17377(.a(new_n17570), .b(new_n17307), .O(new_n17571));
  inv1 g17378(.a(new_n17304), .O(new_n17572));
  nor2 g17379(.a(new_n8170), .b(new_n2660), .O(new_n17573));
  inv1 g17380(.a(new_n17573), .O(new_n17574));
  nor2 g17381(.a(new_n17574), .b(new_n17572), .O(new_n17575));
  nor2 g17382(.a(new_n17575), .b(new_n17571), .O(new_n17576));
  nor2 g17383(.a(new_n17576), .b(new_n17569), .O(new_n17577));
  inv1 g17384(.a(new_n17576), .O(new_n17578));
  nor2 g17385(.a(new_n17578), .b(new_n17568), .O(new_n17579));
  nor2 g17386(.a(new_n17579), .b(new_n17577), .O(new_n17580));
  nor2 g17387(.a(new_n17580), .b(new_n17567), .O(new_n17581));
  inv1 g17388(.a(new_n17567), .O(new_n17582));
  inv1 g17389(.a(new_n17580), .O(new_n17583));
  nor2 g17390(.a(new_n17583), .b(new_n17582), .O(new_n17584));
  nor2 g17391(.a(new_n17584), .b(new_n17581), .O(new_n17585));
  nor2 g17392(.a(new_n17585), .b(new_n17557), .O(new_n17586));
  inv1 g17393(.a(new_n17585), .O(new_n17587));
  nor2 g17394(.a(new_n17587), .b(new_n17556), .O(new_n17588));
  nor2 g17395(.a(new_n17588), .b(new_n17586), .O(new_n17589));
  nor2 g17396(.a(new_n17589), .b(new_n17544), .O(new_n17590));
  inv1 g17397(.a(new_n17544), .O(new_n17591));
  inv1 g17398(.a(new_n17589), .O(new_n17592));
  nor2 g17399(.a(new_n17592), .b(new_n17591), .O(new_n17593));
  nor2 g17400(.a(new_n17593), .b(new_n17590), .O(new_n17594));
  inv1 g17401(.a(new_n17594), .O(new_n17595));
  nor2 g17402(.a(new_n17595), .b(new_n17492), .O(new_n17596));
  inv1 g17403(.a(new_n17492), .O(new_n17597));
  nor2 g17404(.a(new_n17594), .b(new_n17597), .O(new_n17598));
  nor2 g17405(.a(new_n17598), .b(new_n17596), .O(new_n17599));
  inv1 g17406(.a(new_n17599), .O(new_n17600));
  nor2 g17407(.a(new_n17600), .b(new_n17491), .O(new_n17601));
  inv1 g17408(.a(new_n17491), .O(new_n17602));
  nor2 g17409(.a(new_n17599), .b(new_n17602), .O(new_n17603));
  nor2 g17410(.a(new_n17603), .b(new_n17601), .O(new_n17604));
  inv1 g17411(.a(new_n17604), .O(new_n17605));
  nor2 g17412(.a(new_n17605), .b(new_n17490), .O(new_n17606));
  inv1 g17413(.a(new_n17490), .O(new_n17607));
  nor2 g17414(.a(new_n17604), .b(new_n17607), .O(new_n17608));
  nor2 g17415(.a(new_n17608), .b(new_n17606), .O(new_n17609));
  inv1 g17416(.a(new_n17609), .O(new_n17610));
  nor2 g17417(.a(new_n17322), .b(new_n17268), .O(new_n17611));
  inv1 g17418(.a(new_n17611), .O(new_n17612));
  nor2 g17419(.a(new_n17238), .b(new_n17231), .O(new_n17613));
  nor2 g17420(.a(new_n17381), .b(new_n17373), .O(new_n17614));
  nor2 g17421(.a(new_n17614), .b(new_n17613), .O(new_n17615));
  inv1 g17422(.a(new_n17613), .O(new_n17616));
  inv1 g17423(.a(new_n17614), .O(new_n17617));
  nor2 g17424(.a(new_n17617), .b(new_n17616), .O(new_n17618));
  nor2 g17425(.a(new_n17618), .b(new_n17615), .O(new_n17619));
  nor2 g17426(.a(new_n17313), .b(new_n17305), .O(new_n17620));
  nor2 g17427(.a(new_n17620), .b(new_n17619), .O(new_n17621));
  inv1 g17428(.a(new_n17619), .O(new_n17622));
  inv1 g17429(.a(new_n17620), .O(new_n17623));
  nor2 g17430(.a(new_n17623), .b(new_n17622), .O(new_n17624));
  nor2 g17431(.a(new_n17624), .b(new_n17621), .O(new_n17625));
  inv1 g17432(.a(new_n17625), .O(new_n17626));
  nor2 g17433(.a(new_n17250), .b(new_n17242), .O(new_n17627));
  nor2 g17434(.a(new_n17279), .b(new_n17273), .O(new_n17628));
  nor2 g17435(.a(new_n17628), .b(new_n17627), .O(new_n17629));
  inv1 g17436(.a(new_n17627), .O(new_n17630));
  inv1 g17437(.a(new_n17628), .O(new_n17631));
  nor2 g17438(.a(new_n17631), .b(new_n17630), .O(new_n17632));
  nor2 g17439(.a(new_n17632), .b(new_n17629), .O(new_n17633));
  nor2 g17440(.a(new_n17294), .b(new_n17286), .O(new_n17634));
  nor2 g17441(.a(new_n17634), .b(new_n17633), .O(new_n17635));
  inv1 g17442(.a(new_n17633), .O(new_n17636));
  inv1 g17443(.a(new_n17634), .O(new_n17637));
  nor2 g17444(.a(new_n17637), .b(new_n17636), .O(new_n17638));
  nor2 g17445(.a(new_n17638), .b(new_n17635), .O(new_n17639));
  nor2 g17446(.a(new_n17315), .b(new_n17296), .O(new_n17640));
  inv1 g17447(.a(new_n17640), .O(new_n17641));
  nor2 g17448(.a(new_n17641), .b(new_n17639), .O(new_n17642));
  inv1 g17449(.a(new_n17639), .O(new_n17643));
  nor2 g17450(.a(new_n17640), .b(new_n17643), .O(new_n17644));
  nor2 g17451(.a(new_n17644), .b(new_n17642), .O(new_n17645));
  inv1 g17452(.a(new_n17645), .O(new_n17646));
  nor2 g17453(.a(new_n17646), .b(new_n17626), .O(new_n17647));
  nor2 g17454(.a(new_n17645), .b(new_n17625), .O(new_n17648));
  nor2 g17455(.a(new_n17648), .b(new_n17647), .O(new_n17649));
  nor2 g17456(.a(new_n17649), .b(new_n17612), .O(new_n17650));
  inv1 g17457(.a(new_n17649), .O(new_n17651));
  nor2 g17458(.a(new_n17651), .b(new_n17611), .O(new_n17652));
  nor2 g17459(.a(new_n17652), .b(new_n17650), .O(new_n17653));
  inv1 g17460(.a(new_n17653), .O(new_n17654));
  nor2 g17461(.a(new_n17264), .b(new_n17257), .O(new_n17655));
  inv1 g17462(.a(new_n17655), .O(new_n17656));
  nor2 g17463(.a(new_n17383), .b(new_n17367), .O(new_n17657));
  inv1 g17464(.a(new_n17657), .O(new_n17658));
  nor2 g17465(.a(new_n17658), .b(new_n17656), .O(new_n17659));
  nor2 g17466(.a(new_n17657), .b(new_n17655), .O(new_n17660));
  nor2 g17467(.a(new_n17660), .b(new_n17659), .O(new_n17661));
  inv1 g17468(.a(new_n17661), .O(new_n17662));
  nor2 g17469(.a(new_n17255), .b(new_n4954), .O(new_n17663));
  inv1 g17470(.a(new_n17663), .O(new_n17664));
  nor2 g17471(.a(new_n17664), .b(new_n15607), .O(new_n17665));
  nor2 g17472(.a(new_n17663), .b(new_n15606), .O(new_n17666));
  nor2 g17473(.a(new_n17666), .b(new_n17665), .O(new_n17667));
  nor2 g17474(.a(new_n17441), .b(new_n17433), .O(new_n17668));
  nor2 g17475(.a(new_n17668), .b(new_n17667), .O(new_n17669));
  inv1 g17476(.a(new_n17667), .O(new_n17670));
  inv1 g17477(.a(new_n17668), .O(new_n17671));
  nor2 g17478(.a(new_n17671), .b(new_n17670), .O(new_n17672));
  nor2 g17479(.a(new_n17672), .b(new_n17669), .O(new_n17673));
  inv1 g17480(.a(new_n17673), .O(new_n17674));
  nor2 g17481(.a(new_n17674), .b(new_n17662), .O(new_n17675));
  nor2 g17482(.a(new_n17673), .b(new_n17661), .O(new_n17676));
  nor2 g17483(.a(new_n17676), .b(new_n17675), .O(new_n17677));
  inv1 g17484(.a(new_n17677), .O(new_n17678));
  nor2 g17485(.a(new_n17678), .b(new_n17654), .O(new_n17679));
  nor2 g17486(.a(new_n17677), .b(new_n17653), .O(new_n17680));
  nor2 g17487(.a(new_n17680), .b(new_n17679), .O(new_n17681));
  inv1 g17488(.a(new_n17681), .O(new_n17682));
  nor2 g17489(.a(new_n17330), .b(new_n17325), .O(new_n17683));
  nor2 g17490(.a(new_n17407), .b(new_n17401), .O(new_n17684));
  inv1 g17491(.a(new_n17684), .O(new_n17685));
  nor2 g17492(.a(new_n17353), .b(new_n17347), .O(new_n17686));
  nor2 g17493(.a(new_n8946), .b(new_n2184), .O(new_n17687));
  nor2 g17494(.a(new_n9658), .b(new_n1903), .O(new_n17688));
  nor2 g17495(.a(new_n17688), .b(new_n17687), .O(new_n17689));
  nor2 g17496(.a(new_n9658), .b(new_n2184), .O(new_n17690));
  inv1 g17497(.a(new_n17690), .O(new_n17691));
  nor2 g17498(.a(new_n17691), .b(new_n17067), .O(new_n17692));
  nor2 g17499(.a(new_n17692), .b(new_n17689), .O(new_n17693));
  nor2 g17500(.a(new_n17693), .b(new_n8748), .O(new_n17694));
  inv1 g17501(.a(new_n17693), .O(new_n17695));
  nor2 g17502(.a(new_n17695), .b(new_n8747), .O(new_n17696));
  nor2 g17503(.a(new_n17696), .b(new_n17694), .O(new_n17697));
  nor2 g17504(.a(new_n17697), .b(new_n17686), .O(new_n17698));
  inv1 g17505(.a(new_n17686), .O(new_n17699));
  inv1 g17506(.a(new_n17697), .O(new_n17700));
  nor2 g17507(.a(new_n17700), .b(new_n17699), .O(new_n17701));
  nor2 g17508(.a(new_n17701), .b(new_n17698), .O(new_n17702));
  nor2 g17509(.a(new_n17702), .b(new_n17685), .O(new_n17703));
  inv1 g17510(.a(new_n17702), .O(new_n17704));
  nor2 g17511(.a(new_n17704), .b(new_n17684), .O(new_n17705));
  nor2 g17512(.a(new_n17705), .b(new_n17703), .O(new_n17706));
  inv1 g17513(.a(new_n17706), .O(new_n17707));
  nor2 g17514(.a(new_n17418), .b(new_n17415), .O(new_n17708));
  nor2 g17515(.a(new_n17388), .b(new_n17357), .O(new_n17709));
  nor2 g17516(.a(new_n17709), .b(new_n17708), .O(new_n17710));
  inv1 g17517(.a(new_n17708), .O(new_n17711));
  inv1 g17518(.a(new_n17709), .O(new_n17712));
  nor2 g17519(.a(new_n17712), .b(new_n17711), .O(new_n17713));
  nor2 g17520(.a(new_n17713), .b(new_n17710), .O(new_n17714));
  inv1 g17521(.a(new_n17714), .O(new_n17715));
  nor2 g17522(.a(new_n17715), .b(new_n17707), .O(new_n17716));
  nor2 g17523(.a(new_n17714), .b(new_n17706), .O(new_n17717));
  nor2 g17524(.a(new_n17717), .b(new_n17716), .O(new_n17718));
  inv1 g17525(.a(new_n17718), .O(new_n17719));
  nor2 g17526(.a(new_n17719), .b(new_n17683), .O(new_n17720));
  inv1 g17527(.a(new_n17683), .O(new_n17721));
  nor2 g17528(.a(new_n17718), .b(new_n17721), .O(new_n17722));
  nor2 g17529(.a(new_n17722), .b(new_n17720), .O(new_n17723));
  inv1 g17530(.a(new_n17723), .O(new_n17724));
  nor2 g17531(.a(new_n17724), .b(new_n17682), .O(new_n17725));
  nor2 g17532(.a(new_n17723), .b(new_n17681), .O(new_n17726));
  nor2 g17533(.a(new_n17726), .b(new_n17725), .O(new_n17727));
  inv1 g17534(.a(new_n17727), .O(new_n17728));
  nor2 g17535(.a(new_n17728), .b(new_n17610), .O(new_n17729));
  nor2 g17536(.a(new_n17727), .b(new_n17609), .O(new_n17730));
  nor2 g17537(.a(new_n17730), .b(new_n17729), .O(new_n17731));
  inv1 g17538(.a(new_n17731), .O(new_n17732));
  nor2 g17539(.a(new_n17732), .b(new_n17489), .O(new_n17733));
  inv1 g17540(.a(new_n17489), .O(new_n17734));
  nor2 g17541(.a(new_n17731), .b(new_n17734), .O(new_n17735));
  nor2 g17542(.a(new_n17735), .b(new_n17733), .O(new_n17736));
  nor2 g17543(.a(new_n17484), .b(new_n17480), .O(new_n17737));
  inv1 g17544(.a(new_n17737), .O(new_n17738));
  nor2 g17545(.a(new_n17738), .b(new_n17736), .O(new_n17739));
  inv1 g17546(.a(new_n17736), .O(new_n17740));
  nor2 g17547(.a(new_n17737), .b(new_n17740), .O(new_n17741));
  nor2 g17548(.a(new_n17741), .b(new_n17739), .O(new_n17742));
  inv1 g17549(.a(new_n17742), .O(\asquared[83] ));
  nor2 g17550(.a(new_n17729), .b(new_n17606), .O(new_n17744));
  nor2 g17551(.a(new_n17725), .b(new_n17720), .O(new_n17745));
  nor2 g17552(.a(new_n17679), .b(new_n17652), .O(new_n17746));
  nor2 g17553(.a(new_n17716), .b(new_n17710), .O(new_n17747));
  nor2 g17554(.a(new_n17705), .b(new_n17698), .O(new_n17748));
  inv1 g17555(.a(new_n17748), .O(new_n17749));
  nor2 g17556(.a(new_n7294), .b(new_n3231), .O(new_n17750));
  inv1 g17557(.a(new_n17750), .O(new_n17751));
  nor2 g17558(.a(new_n6893), .b(new_n3722), .O(new_n17752));
  nor2 g17559(.a(new_n17752), .b(new_n17513), .O(new_n17753));
  nor2 g17560(.a(new_n6958), .b(new_n3722), .O(new_n17754));
  inv1 g17561(.a(new_n17754), .O(new_n17755));
  nor2 g17562(.a(new_n17755), .b(new_n17233), .O(new_n17756));
  nor2 g17563(.a(new_n17756), .b(new_n17753), .O(new_n17757));
  nor2 g17564(.a(new_n17757), .b(new_n17751), .O(new_n17758));
  inv1 g17565(.a(new_n17757), .O(new_n17759));
  nor2 g17566(.a(new_n17759), .b(new_n17750), .O(new_n17760));
  nor2 g17567(.a(new_n17760), .b(new_n17758), .O(new_n17761));
  inv1 g17568(.a(new_n17761), .O(new_n17762));
  nor2 g17569(.a(new_n8476), .b(new_n2506), .O(new_n17763));
  inv1 g17570(.a(new_n17763), .O(new_n17764));
  nor2 g17571(.a(new_n5393), .b(new_n4682), .O(new_n17765));
  nor2 g17572(.a(new_n17765), .b(new_n17560), .O(new_n17766));
  nor2 g17573(.a(new_n5796), .b(new_n4682), .O(new_n17767));
  inv1 g17574(.a(new_n17767), .O(new_n17768));
  nor2 g17575(.a(new_n17768), .b(new_n17436), .O(new_n17769));
  nor2 g17576(.a(new_n17769), .b(new_n17766), .O(new_n17770));
  nor2 g17577(.a(new_n17770), .b(new_n17764), .O(new_n17771));
  inv1 g17578(.a(new_n17770), .O(new_n17772));
  nor2 g17579(.a(new_n17772), .b(new_n17763), .O(new_n17773));
  nor2 g17580(.a(new_n17773), .b(new_n17771), .O(new_n17774));
  nor2 g17581(.a(new_n11186), .b(new_n1425), .O(new_n17775));
  inv1 g17582(.a(new_n17775), .O(new_n17776));
  nor2 g17583(.a(new_n5178), .b(\a[41] ), .O(new_n17777));
  nor2 g17584(.a(new_n17777), .b(new_n17776), .O(new_n17778));
  inv1 g17585(.a(new_n17777), .O(new_n17779));
  nor2 g17586(.a(new_n17779), .b(new_n17775), .O(new_n17780));
  nor2 g17587(.a(new_n17780), .b(new_n17778), .O(new_n17781));
  nor2 g17588(.a(new_n17781), .b(new_n17774), .O(new_n17782));
  inv1 g17589(.a(new_n17774), .O(new_n17783));
  inv1 g17590(.a(new_n17781), .O(new_n17784));
  nor2 g17591(.a(new_n17784), .b(new_n17783), .O(new_n17785));
  nor2 g17592(.a(new_n17785), .b(new_n17782), .O(new_n17786));
  nor2 g17593(.a(new_n17786), .b(new_n17762), .O(new_n17787));
  inv1 g17594(.a(new_n17786), .O(new_n17788));
  nor2 g17595(.a(new_n17788), .b(new_n17761), .O(new_n17789));
  nor2 g17596(.a(new_n17789), .b(new_n17787), .O(new_n17790));
  nor2 g17597(.a(new_n17790), .b(new_n17749), .O(new_n17791));
  inv1 g17598(.a(new_n17790), .O(new_n17792));
  nor2 g17599(.a(new_n17792), .b(new_n17748), .O(new_n17793));
  nor2 g17600(.a(new_n17793), .b(new_n17791), .O(new_n17794));
  nor2 g17601(.a(new_n11596), .b(new_n1297), .O(new_n17795));
  nor2 g17602(.a(new_n10895), .b(new_n1493), .O(new_n17796));
  nor2 g17603(.a(new_n17796), .b(new_n17795), .O(new_n17797));
  inv1 g17604(.a(new_n17271), .O(new_n17798));
  nor2 g17605(.a(new_n11596), .b(new_n1493), .O(new_n17799));
  inv1 g17606(.a(new_n17799), .O(new_n17800));
  nor2 g17607(.a(new_n17800), .b(new_n17798), .O(new_n17801));
  nor2 g17608(.a(new_n17801), .b(new_n17797), .O(new_n17802));
  nor2 g17609(.a(new_n17802), .b(new_n16714), .O(new_n17803));
  inv1 g17610(.a(new_n17802), .O(new_n17804));
  nor2 g17611(.a(new_n17804), .b(new_n16713), .O(new_n17805));
  nor2 g17612(.a(new_n17805), .b(new_n17803), .O(new_n17806));
  inv1 g17613(.a(new_n17806), .O(new_n17807));
  nor2 g17614(.a(new_n7537), .b(new_n3057), .O(new_n17808));
  nor2 g17615(.a(new_n17808), .b(new_n15680), .O(new_n17809));
  nor2 g17616(.a(new_n9658), .b(new_n3057), .O(new_n17810));
  inv1 g17617(.a(new_n17810), .O(new_n17811));
  nor2 g17618(.a(new_n17811), .b(new_n16132), .O(new_n17812));
  nor2 g17619(.a(new_n17812), .b(new_n17809), .O(new_n17813));
  inv1 g17620(.a(new_n17813), .O(new_n17814));
  nor2 g17621(.a(new_n17814), .b(new_n17244), .O(new_n17815));
  nor2 g17622(.a(new_n17813), .b(new_n17245), .O(new_n17816));
  nor2 g17623(.a(new_n17816), .b(new_n17815), .O(new_n17817));
  nor2 g17624(.a(new_n6570), .b(new_n3870), .O(new_n17818));
  inv1 g17625(.a(new_n17818), .O(new_n17819));
  nor2 g17626(.a(new_n5971), .b(new_n4366), .O(new_n17820));
  nor2 g17627(.a(new_n17820), .b(new_n17549), .O(new_n17821));
  nor2 g17628(.a(new_n6274), .b(new_n4366), .O(new_n17822));
  inv1 g17629(.a(new_n17822), .O(new_n17823));
  nor2 g17630(.a(new_n17823), .b(new_n17289), .O(new_n17824));
  nor2 g17631(.a(new_n17824), .b(new_n17821), .O(new_n17825));
  nor2 g17632(.a(new_n17825), .b(new_n17819), .O(new_n17826));
  inv1 g17633(.a(new_n17825), .O(new_n17827));
  nor2 g17634(.a(new_n17827), .b(new_n17818), .O(new_n17828));
  nor2 g17635(.a(new_n17828), .b(new_n17826), .O(new_n17829));
  nor2 g17636(.a(new_n17829), .b(new_n17817), .O(new_n17830));
  inv1 g17637(.a(new_n17817), .O(new_n17831));
  inv1 g17638(.a(new_n17829), .O(new_n17832));
  nor2 g17639(.a(new_n17832), .b(new_n17831), .O(new_n17833));
  nor2 g17640(.a(new_n17833), .b(new_n17830), .O(new_n17834));
  nor2 g17641(.a(new_n17834), .b(new_n17807), .O(new_n17835));
  inv1 g17642(.a(new_n17834), .O(new_n17836));
  nor2 g17643(.a(new_n17836), .b(new_n17806), .O(new_n17837));
  nor2 g17644(.a(new_n17837), .b(new_n17835), .O(new_n17838));
  nor2 g17645(.a(new_n17838), .b(new_n17794), .O(new_n17839));
  inv1 g17646(.a(new_n17794), .O(new_n17840));
  inv1 g17647(.a(new_n17838), .O(new_n17841));
  nor2 g17648(.a(new_n17841), .b(new_n17840), .O(new_n17842));
  nor2 g17649(.a(new_n17842), .b(new_n17839), .O(new_n17843));
  inv1 g17650(.a(new_n17843), .O(new_n17844));
  nor2 g17651(.a(new_n17844), .b(new_n17747), .O(new_n17845));
  inv1 g17652(.a(new_n17747), .O(new_n17846));
  nor2 g17653(.a(new_n17843), .b(new_n17846), .O(new_n17847));
  nor2 g17654(.a(new_n17847), .b(new_n17845), .O(new_n17848));
  inv1 g17655(.a(new_n17848), .O(new_n17849));
  nor2 g17656(.a(new_n17849), .b(new_n17746), .O(new_n17850));
  inv1 g17657(.a(new_n17746), .O(new_n17851));
  nor2 g17658(.a(new_n17848), .b(new_n17851), .O(new_n17852));
  nor2 g17659(.a(new_n17852), .b(new_n17850), .O(new_n17853));
  inv1 g17660(.a(new_n17853), .O(new_n17854));
  nor2 g17661(.a(new_n17854), .b(new_n17745), .O(new_n17855));
  inv1 g17662(.a(new_n17745), .O(new_n17856));
  nor2 g17663(.a(new_n17853), .b(new_n17856), .O(new_n17857));
  nor2 g17664(.a(new_n17857), .b(new_n17855), .O(new_n17858));
  inv1 g17665(.a(new_n17858), .O(new_n17859));
  nor2 g17666(.a(new_n17601), .b(new_n17596), .O(new_n17860));
  nor2 g17667(.a(new_n17624), .b(new_n17618), .O(new_n17861));
  inv1 g17668(.a(new_n17861), .O(new_n17862));
  nor2 g17669(.a(new_n17638), .b(new_n17632), .O(new_n17863));
  inv1 g17670(.a(new_n17863), .O(new_n17864));
  nor2 g17671(.a(new_n17864), .b(new_n17862), .O(new_n17865));
  nor2 g17672(.a(new_n17863), .b(new_n17861), .O(new_n17866));
  nor2 g17673(.a(new_n17866), .b(new_n17865), .O(new_n17867));
  nor2 g17674(.a(new_n17539), .b(new_n17532), .O(new_n17868));
  inv1 g17675(.a(new_n17868), .O(new_n17869));
  nor2 g17676(.a(new_n17869), .b(new_n17867), .O(new_n17870));
  inv1 g17677(.a(new_n17867), .O(new_n17871));
  nor2 g17678(.a(new_n17868), .b(new_n17871), .O(new_n17872));
  nor2 g17679(.a(new_n17872), .b(new_n17870), .O(new_n17873));
  inv1 g17680(.a(new_n17873), .O(new_n17874));
  nor2 g17681(.a(new_n17672), .b(new_n17665), .O(new_n17875));
  inv1 g17682(.a(new_n17875), .O(new_n17876));
  nor2 g17683(.a(new_n8026), .b(new_n2826), .O(new_n17877));
  inv1 g17684(.a(new_n17877), .O(new_n17878));
  nor2 g17685(.a(new_n8946), .b(new_n2433), .O(new_n17879));
  nor2 g17686(.a(new_n17879), .b(new_n17573), .O(new_n17880));
  nor2 g17687(.a(new_n8946), .b(new_n2660), .O(new_n17881));
  inv1 g17688(.a(new_n17881), .O(new_n17882));
  nor2 g17689(.a(new_n17882), .b(new_n17047), .O(new_n17883));
  nor2 g17690(.a(new_n17883), .b(new_n17880), .O(new_n17884));
  nor2 g17691(.a(new_n17884), .b(new_n17878), .O(new_n17885));
  inv1 g17692(.a(new_n17884), .O(new_n17886));
  nor2 g17693(.a(new_n17886), .b(new_n17877), .O(new_n17887));
  nor2 g17694(.a(new_n17887), .b(new_n17885), .O(new_n17888));
  nor2 g17695(.a(new_n10468), .b(new_n1647), .O(new_n17889));
  nor2 g17696(.a(new_n17889), .b(new_n17501), .O(new_n17890));
  inv1 g17697(.a(new_n17498), .O(new_n17891));
  nor2 g17698(.a(new_n10468), .b(new_n1736), .O(new_n17892));
  inv1 g17699(.a(new_n17892), .O(new_n17893));
  nor2 g17700(.a(new_n17893), .b(new_n17891), .O(new_n17894));
  nor2 g17701(.a(new_n17894), .b(new_n17890), .O(new_n17895));
  inv1 g17702(.a(new_n17895), .O(new_n17896));
  nor2 g17703(.a(new_n17579), .b(new_n17571), .O(new_n17897));
  inv1 g17704(.a(new_n17897), .O(new_n17898));
  nor2 g17705(.a(new_n17898), .b(new_n17896), .O(new_n17899));
  nor2 g17706(.a(new_n17897), .b(new_n17895), .O(new_n17900));
  nor2 g17707(.a(new_n17900), .b(new_n17899), .O(new_n17901));
  inv1 g17708(.a(new_n17901), .O(new_n17902));
  nor2 g17709(.a(new_n17902), .b(new_n17888), .O(new_n17903));
  inv1 g17710(.a(new_n17888), .O(new_n17904));
  nor2 g17711(.a(new_n17901), .b(new_n17904), .O(new_n17905));
  nor2 g17712(.a(new_n17905), .b(new_n17903), .O(new_n17906));
  nor2 g17713(.a(new_n17906), .b(new_n17876), .O(new_n17907));
  inv1 g17714(.a(new_n17906), .O(new_n17908));
  nor2 g17715(.a(new_n17908), .b(new_n17875), .O(new_n17909));
  nor2 g17716(.a(new_n17909), .b(new_n17907), .O(new_n17910));
  inv1 g17717(.a(new_n17910), .O(new_n17911));
  nor2 g17718(.a(new_n17675), .b(new_n17660), .O(new_n17912));
  nor2 g17719(.a(new_n17912), .b(new_n17911), .O(new_n17913));
  inv1 g17720(.a(new_n17912), .O(new_n17914));
  nor2 g17721(.a(new_n17914), .b(new_n17910), .O(new_n17915));
  nor2 g17722(.a(new_n17915), .b(new_n17913), .O(new_n17916));
  inv1 g17723(.a(new_n17916), .O(new_n17917));
  nor2 g17724(.a(new_n17917), .b(new_n17874), .O(new_n17918));
  nor2 g17725(.a(new_n17916), .b(new_n17873), .O(new_n17919));
  nor2 g17726(.a(new_n17919), .b(new_n17918), .O(new_n17920));
  inv1 g17727(.a(new_n17920), .O(new_n17921));
  nor2 g17728(.a(new_n17921), .b(new_n17860), .O(new_n17922));
  inv1 g17729(.a(new_n17860), .O(new_n17923));
  nor2 g17730(.a(new_n17920), .b(new_n17923), .O(new_n17924));
  nor2 g17731(.a(new_n17924), .b(new_n17922), .O(new_n17925));
  nor2 g17732(.a(new_n17507), .b(new_n17499), .O(new_n17926));
  nor2 g17733(.a(new_n17555), .b(new_n17548), .O(new_n17927));
  nor2 g17734(.a(new_n17927), .b(new_n17926), .O(new_n17928));
  inv1 g17735(.a(new_n17926), .O(new_n17929));
  inv1 g17736(.a(new_n17927), .O(new_n17930));
  nor2 g17737(.a(new_n17930), .b(new_n17929), .O(new_n17931));
  nor2 g17738(.a(new_n17931), .b(new_n17928), .O(new_n17932));
  nor2 g17739(.a(new_n17565), .b(new_n17559), .O(new_n17933));
  nor2 g17740(.a(new_n17933), .b(new_n17932), .O(new_n17934));
  inv1 g17741(.a(new_n17932), .O(new_n17935));
  inv1 g17742(.a(new_n17933), .O(new_n17936));
  nor2 g17743(.a(new_n17936), .b(new_n17935), .O(new_n17937));
  nor2 g17744(.a(new_n17937), .b(new_n17934), .O(new_n17938));
  inv1 g17745(.a(new_n17938), .O(new_n17939));
  nor2 g17746(.a(new_n17530), .b(new_n17524), .O(new_n17940));
  nor2 g17747(.a(new_n17519), .b(new_n17511), .O(new_n17941));
  nor2 g17748(.a(new_n17941), .b(new_n17940), .O(new_n17942));
  inv1 g17749(.a(new_n17940), .O(new_n17943));
  inv1 g17750(.a(new_n17941), .O(new_n17944));
  nor2 g17751(.a(new_n17944), .b(new_n17943), .O(new_n17945));
  nor2 g17752(.a(new_n17945), .b(new_n17942), .O(new_n17946));
  nor2 g17753(.a(new_n17696), .b(new_n17689), .O(new_n17947));
  nor2 g17754(.a(new_n17947), .b(new_n17946), .O(new_n17948));
  inv1 g17755(.a(new_n17946), .O(new_n17949));
  inv1 g17756(.a(new_n17947), .O(new_n17950));
  nor2 g17757(.a(new_n17950), .b(new_n17949), .O(new_n17951));
  nor2 g17758(.a(new_n17951), .b(new_n17948), .O(new_n17952));
  nor2 g17759(.a(new_n17588), .b(new_n17581), .O(new_n17953));
  inv1 g17760(.a(new_n17953), .O(new_n17954));
  nor2 g17761(.a(new_n17954), .b(new_n17952), .O(new_n17955));
  inv1 g17762(.a(new_n17952), .O(new_n17956));
  nor2 g17763(.a(new_n17953), .b(new_n17956), .O(new_n17957));
  nor2 g17764(.a(new_n17957), .b(new_n17955), .O(new_n17958));
  inv1 g17765(.a(new_n17958), .O(new_n17959));
  nor2 g17766(.a(new_n17959), .b(new_n17939), .O(new_n17960));
  nor2 g17767(.a(new_n17958), .b(new_n17938), .O(new_n17961));
  nor2 g17768(.a(new_n17961), .b(new_n17960), .O(new_n17962));
  inv1 g17769(.a(new_n17962), .O(new_n17963));
  nor2 g17770(.a(new_n17593), .b(new_n17543), .O(new_n17964));
  nor2 g17771(.a(new_n17647), .b(new_n17644), .O(new_n17965));
  nor2 g17772(.a(new_n17965), .b(new_n17964), .O(new_n17966));
  inv1 g17773(.a(new_n17964), .O(new_n17967));
  inv1 g17774(.a(new_n17965), .O(new_n17968));
  nor2 g17775(.a(new_n17968), .b(new_n17967), .O(new_n17969));
  nor2 g17776(.a(new_n17969), .b(new_n17966), .O(new_n17970));
  inv1 g17777(.a(new_n17970), .O(new_n17971));
  nor2 g17778(.a(new_n17971), .b(new_n17963), .O(new_n17972));
  nor2 g17779(.a(new_n17970), .b(new_n17962), .O(new_n17973));
  nor2 g17780(.a(new_n17973), .b(new_n17972), .O(new_n17974));
  inv1 g17781(.a(new_n17974), .O(new_n17975));
  nor2 g17782(.a(new_n17975), .b(new_n17925), .O(new_n17976));
  inv1 g17783(.a(new_n17925), .O(new_n17977));
  nor2 g17784(.a(new_n17974), .b(new_n17977), .O(new_n17978));
  nor2 g17785(.a(new_n17978), .b(new_n17976), .O(new_n17979));
  nor2 g17786(.a(new_n17979), .b(new_n17859), .O(new_n17980));
  inv1 g17787(.a(new_n17979), .O(new_n17981));
  nor2 g17788(.a(new_n17981), .b(new_n17858), .O(new_n17982));
  nor2 g17789(.a(new_n17982), .b(new_n17980), .O(new_n17983));
  inv1 g17790(.a(new_n17983), .O(new_n17984));
  nor2 g17791(.a(new_n17984), .b(new_n17744), .O(new_n17985));
  inv1 g17792(.a(new_n17744), .O(new_n17986));
  nor2 g17793(.a(new_n17983), .b(new_n17986), .O(new_n17987));
  nor2 g17794(.a(new_n17987), .b(new_n17985), .O(new_n17988));
  inv1 g17795(.a(new_n17988), .O(new_n17989));
  nor2 g17796(.a(new_n17741), .b(new_n17735), .O(new_n17990));
  nor2 g17797(.a(new_n17990), .b(new_n17989), .O(new_n17991));
  inv1 g17798(.a(new_n17990), .O(new_n17992));
  nor2 g17799(.a(new_n17992), .b(new_n17988), .O(new_n17993));
  nor2 g17800(.a(new_n17993), .b(new_n17991), .O(new_n17994));
  inv1 g17801(.a(new_n17994), .O(\asquared[84] ));
  nor2 g17802(.a(new_n17850), .b(new_n17845), .O(new_n17996));
  inv1 g17803(.a(new_n17996), .O(new_n17997));
  nor2 g17804(.a(new_n17972), .b(new_n17966), .O(new_n17998));
  inv1 g17805(.a(new_n17998), .O(new_n17999));
  nor2 g17806(.a(new_n17999), .b(new_n17997), .O(new_n18000));
  nor2 g17807(.a(new_n17998), .b(new_n17996), .O(new_n18001));
  nor2 g17808(.a(new_n18001), .b(new_n18000), .O(new_n18002));
  inv1 g17809(.a(new_n18002), .O(new_n18003));
  nor2 g17810(.a(new_n17780), .b(new_n5178), .O(new_n18004));
  nor2 g17811(.a(new_n17773), .b(new_n17766), .O(new_n18005));
  nor2 g17812(.a(new_n18005), .b(new_n18004), .O(new_n18006));
  inv1 g17813(.a(new_n18004), .O(new_n18007));
  inv1 g17814(.a(new_n18005), .O(new_n18008));
  nor2 g17815(.a(new_n18008), .b(new_n18007), .O(new_n18009));
  nor2 g17816(.a(new_n18009), .b(new_n18006), .O(new_n18010));
  nor2 g17817(.a(new_n17887), .b(new_n17880), .O(new_n18011));
  nor2 g17818(.a(new_n18011), .b(new_n18010), .O(new_n18012));
  inv1 g17819(.a(new_n18010), .O(new_n18013));
  inv1 g17820(.a(new_n18011), .O(new_n18014));
  nor2 g17821(.a(new_n18014), .b(new_n18013), .O(new_n18015));
  nor2 g17822(.a(new_n18015), .b(new_n18012), .O(new_n18016));
  inv1 g17823(.a(new_n18016), .O(new_n18017));
  nor2 g17824(.a(new_n17837), .b(new_n17830), .O(new_n18018));
  inv1 g17825(.a(new_n18018), .O(new_n18019));
  nor2 g17826(.a(new_n17789), .b(new_n17782), .O(new_n18020));
  inv1 g17827(.a(new_n18020), .O(new_n18021));
  nor2 g17828(.a(new_n18021), .b(new_n18019), .O(new_n18022));
  nor2 g17829(.a(new_n18020), .b(new_n18018), .O(new_n18023));
  nor2 g17830(.a(new_n18023), .b(new_n18022), .O(new_n18024));
  inv1 g17831(.a(new_n18024), .O(new_n18025));
  nor2 g17832(.a(new_n18025), .b(new_n18017), .O(new_n18026));
  nor2 g17833(.a(new_n18024), .b(new_n18016), .O(new_n18027));
  nor2 g17834(.a(new_n18027), .b(new_n18026), .O(new_n18028));
  inv1 g17835(.a(new_n18028), .O(new_n18029));
  nor2 g17836(.a(new_n17842), .b(new_n17793), .O(new_n18030));
  nor2 g17837(.a(new_n17960), .b(new_n17957), .O(new_n18031));
  nor2 g17838(.a(new_n18031), .b(new_n18030), .O(new_n18032));
  inv1 g17839(.a(new_n18030), .O(new_n18033));
  inv1 g17840(.a(new_n18031), .O(new_n18034));
  nor2 g17841(.a(new_n18034), .b(new_n18033), .O(new_n18035));
  nor2 g17842(.a(new_n18035), .b(new_n18032), .O(new_n18036));
  inv1 g17843(.a(new_n18036), .O(new_n18037));
  nor2 g17844(.a(new_n18037), .b(new_n18029), .O(new_n18038));
  nor2 g17845(.a(new_n18036), .b(new_n18028), .O(new_n18039));
  nor2 g17846(.a(new_n18039), .b(new_n18038), .O(new_n18040));
  inv1 g17847(.a(new_n18040), .O(new_n18041));
  nor2 g17848(.a(new_n18041), .b(new_n18003), .O(new_n18042));
  nor2 g17849(.a(new_n18040), .b(new_n18002), .O(new_n18043));
  nor2 g17850(.a(new_n18043), .b(new_n18042), .O(new_n18044));
  inv1 g17851(.a(new_n18044), .O(new_n18045));
  nor2 g17852(.a(new_n17909), .b(new_n17903), .O(new_n18046));
  inv1 g17853(.a(new_n18046), .O(new_n18047));
  nor2 g17854(.a(new_n17899), .b(new_n17894), .O(new_n18048));
  inv1 g17855(.a(new_n18048), .O(new_n18049));
  nor2 g17856(.a(new_n17805), .b(new_n17797), .O(new_n18050));
  nor2 g17857(.a(new_n18050), .b(new_n18049), .O(new_n18051));
  inv1 g17858(.a(new_n18050), .O(new_n18052));
  nor2 g17859(.a(new_n18052), .b(new_n18048), .O(new_n18053));
  nor2 g17860(.a(new_n18053), .b(new_n18051), .O(new_n18054));
  inv1 g17861(.a(new_n18054), .O(new_n18055));
  nor2 g17862(.a(new_n9873), .b(new_n2121), .O(new_n18056));
  inv1 g17863(.a(new_n18056), .O(new_n18057));
  nor2 g17864(.a(new_n8170), .b(new_n2826), .O(new_n18058));
  nor2 g17865(.a(new_n8026), .b(new_n3057), .O(new_n18059));
  nor2 g17866(.a(new_n18059), .b(new_n18058), .O(new_n18060));
  nor2 g17867(.a(new_n8170), .b(new_n3057), .O(new_n18061));
  inv1 g17868(.a(new_n18061), .O(new_n18062));
  nor2 g17869(.a(new_n18062), .b(new_n17878), .O(new_n18063));
  nor2 g17870(.a(new_n18063), .b(new_n18060), .O(new_n18064));
  nor2 g17871(.a(new_n18064), .b(new_n18057), .O(new_n18065));
  inv1 g17872(.a(new_n18064), .O(new_n18066));
  nor2 g17873(.a(new_n18066), .b(new_n18056), .O(new_n18067));
  nor2 g17874(.a(new_n18067), .b(new_n18065), .O(new_n18068));
  nor2 g17875(.a(new_n18068), .b(new_n18055), .O(new_n18069));
  inv1 g17876(.a(new_n18068), .O(new_n18070));
  nor2 g17877(.a(new_n18070), .b(new_n18054), .O(new_n18071));
  nor2 g17878(.a(new_n18071), .b(new_n18069), .O(new_n18072));
  nor2 g17879(.a(new_n18072), .b(new_n18047), .O(new_n18073));
  inv1 g17880(.a(new_n18072), .O(new_n18074));
  nor2 g17881(.a(new_n18074), .b(new_n18046), .O(new_n18075));
  nor2 g17882(.a(new_n18075), .b(new_n18073), .O(new_n18076));
  nor2 g17883(.a(new_n17872), .b(new_n17866), .O(new_n18077));
  inv1 g17884(.a(new_n18077), .O(new_n18078));
  nor2 g17885(.a(new_n18078), .b(new_n18076), .O(new_n18079));
  inv1 g17886(.a(new_n18076), .O(new_n18080));
  nor2 g17887(.a(new_n18077), .b(new_n18080), .O(new_n18081));
  nor2 g17888(.a(new_n18081), .b(new_n18079), .O(new_n18082));
  nor2 g17889(.a(new_n17918), .b(new_n17913), .O(new_n18083));
  inv1 g17890(.a(new_n18083), .O(new_n18084));
  nor2 g17891(.a(new_n18084), .b(new_n18082), .O(new_n18085));
  inv1 g17892(.a(new_n18082), .O(new_n18086));
  nor2 g17893(.a(new_n18083), .b(new_n18086), .O(new_n18087));
  nor2 g17894(.a(new_n18087), .b(new_n18085), .O(new_n18088));
  inv1 g17895(.a(new_n18088), .O(new_n18089));
  nor2 g17896(.a(new_n17760), .b(new_n17753), .O(new_n18090));
  nor2 g17897(.a(new_n17828), .b(new_n17821), .O(new_n18091));
  nor2 g17898(.a(new_n18091), .b(new_n18090), .O(new_n18092));
  inv1 g17899(.a(new_n18090), .O(new_n18093));
  inv1 g17900(.a(new_n18091), .O(new_n18094));
  nor2 g17901(.a(new_n18094), .b(new_n18093), .O(new_n18095));
  nor2 g17902(.a(new_n18095), .b(new_n18092), .O(new_n18096));
  nor2 g17903(.a(new_n17815), .b(new_n17809), .O(new_n18097));
  nor2 g17904(.a(new_n18097), .b(new_n18096), .O(new_n18098));
  inv1 g17905(.a(new_n18096), .O(new_n18099));
  inv1 g17906(.a(new_n18097), .O(new_n18100));
  nor2 g17907(.a(new_n18100), .b(new_n18099), .O(new_n18101));
  nor2 g17908(.a(new_n18101), .b(new_n18098), .O(new_n18102));
  inv1 g17909(.a(new_n18102), .O(new_n18103));
  nor2 g17910(.a(new_n17937), .b(new_n17931), .O(new_n18104));
  inv1 g17911(.a(new_n18104), .O(new_n18105));
  nor2 g17912(.a(new_n17951), .b(new_n17945), .O(new_n18106));
  inv1 g17913(.a(new_n18106), .O(new_n18107));
  nor2 g17914(.a(new_n18107), .b(new_n18105), .O(new_n18108));
  nor2 g17915(.a(new_n18106), .b(new_n18104), .O(new_n18109));
  nor2 g17916(.a(new_n18109), .b(new_n18108), .O(new_n18110));
  inv1 g17917(.a(new_n18110), .O(new_n18111));
  nor2 g17918(.a(new_n18111), .b(new_n18103), .O(new_n18112));
  nor2 g17919(.a(new_n18110), .b(new_n18102), .O(new_n18113));
  nor2 g17920(.a(new_n18113), .b(new_n18112), .O(new_n18114));
  inv1 g17921(.a(new_n18114), .O(new_n18115));
  nor2 g17922(.a(new_n7294), .b(new_n3533), .O(new_n18116));
  inv1 g17923(.a(new_n18116), .O(new_n18117));
  nor2 g17924(.a(new_n6893), .b(new_n3870), .O(new_n18118));
  nor2 g17925(.a(new_n18118), .b(new_n17754), .O(new_n18119));
  inv1 g17926(.a(new_n17752), .O(new_n18120));
  nor2 g17927(.a(new_n6958), .b(new_n3870), .O(new_n18121));
  inv1 g17928(.a(new_n18121), .O(new_n18122));
  nor2 g17929(.a(new_n18122), .b(new_n18120), .O(new_n18123));
  nor2 g17930(.a(new_n18123), .b(new_n18119), .O(new_n18124));
  nor2 g17931(.a(new_n18124), .b(new_n18117), .O(new_n18125));
  inv1 g17932(.a(new_n18124), .O(new_n18126));
  nor2 g17933(.a(new_n18126), .b(new_n18116), .O(new_n18127));
  nor2 g17934(.a(new_n18127), .b(new_n18125), .O(new_n18128));
  inv1 g17935(.a(new_n18128), .O(new_n18129));
  nor2 g17936(.a(new_n11596), .b(new_n1425), .O(new_n18130));
  nor2 g17937(.a(new_n11186), .b(new_n1493), .O(new_n18131));
  nor2 g17938(.a(new_n10895), .b(new_n1647), .O(new_n18132));
  nor2 g17939(.a(new_n18132), .b(new_n18131), .O(new_n18133));
  inv1 g17940(.a(new_n17796), .O(new_n18134));
  nor2 g17941(.a(new_n11186), .b(new_n1647), .O(new_n18135));
  inv1 g17942(.a(new_n18135), .O(new_n18136));
  nor2 g17943(.a(new_n18136), .b(new_n18134), .O(new_n18137));
  nor2 g17944(.a(new_n18137), .b(new_n18133), .O(new_n18138));
  inv1 g17945(.a(new_n18138), .O(new_n18139));
  nor2 g17946(.a(new_n18139), .b(new_n18130), .O(new_n18140));
  inv1 g17947(.a(new_n18130), .O(new_n18141));
  nor2 g17948(.a(new_n18138), .b(new_n18141), .O(new_n18142));
  nor2 g17949(.a(new_n18142), .b(new_n18140), .O(new_n18143));
  nor2 g17950(.a(new_n7537), .b(new_n3231), .O(new_n18144));
  inv1 g17951(.a(new_n18144), .O(new_n18145));
  nor2 g17952(.a(new_n10320), .b(new_n1903), .O(new_n18146));
  nor2 g17953(.a(new_n18146), .b(new_n17892), .O(new_n18147));
  nor2 g17954(.a(new_n10468), .b(new_n1903), .O(new_n18148));
  inv1 g17955(.a(new_n18148), .O(new_n18149));
  nor2 g17956(.a(new_n18149), .b(new_n17502), .O(new_n18150));
  nor2 g17957(.a(new_n18150), .b(new_n18147), .O(new_n18151));
  nor2 g17958(.a(new_n18151), .b(new_n18145), .O(new_n18152));
  inv1 g17959(.a(new_n18151), .O(new_n18153));
  nor2 g17960(.a(new_n18153), .b(new_n18144), .O(new_n18154));
  nor2 g17961(.a(new_n18154), .b(new_n18152), .O(new_n18155));
  nor2 g17962(.a(new_n18155), .b(new_n18143), .O(new_n18156));
  inv1 g17963(.a(new_n18143), .O(new_n18157));
  inv1 g17964(.a(new_n18155), .O(new_n18158));
  nor2 g17965(.a(new_n18158), .b(new_n18157), .O(new_n18159));
  nor2 g17966(.a(new_n18159), .b(new_n18156), .O(new_n18160));
  nor2 g17967(.a(new_n18160), .b(new_n18129), .O(new_n18161));
  inv1 g17968(.a(new_n18160), .O(new_n18162));
  nor2 g17969(.a(new_n18162), .b(new_n18128), .O(new_n18163));
  nor2 g17970(.a(new_n18163), .b(new_n18161), .O(new_n18164));
  inv1 g17971(.a(new_n18164), .O(new_n18165));
  nor2 g17972(.a(new_n6570), .b(new_n4093), .O(new_n18166));
  inv1 g17973(.a(new_n18166), .O(new_n18167));
  nor2 g17974(.a(new_n8476), .b(new_n2660), .O(new_n18168));
  nor2 g17975(.a(new_n18168), .b(new_n17690), .O(new_n18169));
  nor2 g17976(.a(new_n9658), .b(new_n2660), .O(new_n18170));
  inv1 g17977(.a(new_n18170), .O(new_n18171));
  nor2 g17978(.a(new_n18171), .b(new_n17431), .O(new_n18172));
  nor2 g17979(.a(new_n18172), .b(new_n18169), .O(new_n18173));
  nor2 g17980(.a(new_n18173), .b(new_n18167), .O(new_n18174));
  inv1 g17981(.a(new_n18173), .O(new_n18175));
  nor2 g17982(.a(new_n18175), .b(new_n18166), .O(new_n18176));
  nor2 g17983(.a(new_n18176), .b(new_n18174), .O(new_n18177));
  inv1 g17984(.a(new_n18177), .O(new_n18178));
  nor2 g17985(.a(new_n5971), .b(new_n4425), .O(new_n18179));
  inv1 g17986(.a(new_n18179), .O(new_n18180));
  nor2 g17987(.a(new_n5393), .b(new_n4954), .O(new_n18181));
  nor2 g17988(.a(new_n18181), .b(new_n17767), .O(new_n18182));
  inv1 g17989(.a(new_n17765), .O(new_n18183));
  nor2 g17990(.a(new_n5796), .b(new_n4954), .O(new_n18184));
  inv1 g17991(.a(new_n18184), .O(new_n18185));
  nor2 g17992(.a(new_n18185), .b(new_n18183), .O(new_n18186));
  nor2 g17993(.a(new_n18186), .b(new_n18182), .O(new_n18187));
  nor2 g17994(.a(new_n18187), .b(new_n18180), .O(new_n18188));
  inv1 g17995(.a(new_n18187), .O(new_n18189));
  nor2 g17996(.a(new_n18189), .b(new_n18179), .O(new_n18190));
  nor2 g17997(.a(new_n18190), .b(new_n18188), .O(new_n18191));
  nor2 g17998(.a(new_n9156), .b(new_n2433), .O(new_n18192));
  inv1 g17999(.a(new_n18192), .O(new_n18193));
  nor2 g18000(.a(new_n8946), .b(new_n2506), .O(new_n18194));
  nor2 g18001(.a(new_n18194), .b(new_n17822), .O(new_n18195));
  inv1 g18002(.a(new_n18194), .O(new_n18196));
  nor2 g18003(.a(new_n18196), .b(new_n17823), .O(new_n18197));
  nor2 g18004(.a(new_n18197), .b(new_n18195), .O(new_n18198));
  nor2 g18005(.a(new_n18198), .b(new_n18193), .O(new_n18199));
  inv1 g18006(.a(new_n18198), .O(new_n18200));
  nor2 g18007(.a(new_n18200), .b(new_n18192), .O(new_n18201));
  nor2 g18008(.a(new_n18201), .b(new_n18199), .O(new_n18202));
  nor2 g18009(.a(new_n18202), .b(new_n18191), .O(new_n18203));
  inv1 g18010(.a(new_n18191), .O(new_n18204));
  inv1 g18011(.a(new_n18202), .O(new_n18205));
  nor2 g18012(.a(new_n18205), .b(new_n18204), .O(new_n18206));
  nor2 g18013(.a(new_n18206), .b(new_n18203), .O(new_n18207));
  nor2 g18014(.a(new_n18207), .b(new_n18178), .O(new_n18208));
  inv1 g18015(.a(new_n18207), .O(new_n18209));
  nor2 g18016(.a(new_n18209), .b(new_n18177), .O(new_n18210));
  nor2 g18017(.a(new_n18210), .b(new_n18208), .O(new_n18211));
  inv1 g18018(.a(new_n18211), .O(new_n18212));
  nor2 g18019(.a(new_n18212), .b(new_n18165), .O(new_n18213));
  nor2 g18020(.a(new_n18211), .b(new_n18164), .O(new_n18214));
  nor2 g18021(.a(new_n18214), .b(new_n18213), .O(new_n18215));
  inv1 g18022(.a(new_n18215), .O(new_n18216));
  nor2 g18023(.a(new_n18216), .b(new_n18115), .O(new_n18217));
  nor2 g18024(.a(new_n18215), .b(new_n18114), .O(new_n18218));
  nor2 g18025(.a(new_n18218), .b(new_n18217), .O(new_n18219));
  inv1 g18026(.a(new_n18219), .O(new_n18220));
  nor2 g18027(.a(new_n18220), .b(new_n18089), .O(new_n18221));
  nor2 g18028(.a(new_n18219), .b(new_n18088), .O(new_n18222));
  nor2 g18029(.a(new_n18222), .b(new_n18221), .O(new_n18223));
  inv1 g18030(.a(new_n18223), .O(new_n18224));
  nor2 g18031(.a(new_n17978), .b(new_n17924), .O(new_n18225));
  inv1 g18032(.a(new_n18225), .O(new_n18226));
  nor2 g18033(.a(new_n18226), .b(new_n18224), .O(new_n18227));
  nor2 g18034(.a(new_n18225), .b(new_n18223), .O(new_n18228));
  nor2 g18035(.a(new_n18228), .b(new_n18227), .O(new_n18229));
  inv1 g18036(.a(new_n18229), .O(new_n18230));
  nor2 g18037(.a(new_n18230), .b(new_n18045), .O(new_n18231));
  nor2 g18038(.a(new_n18229), .b(new_n18044), .O(new_n18232));
  nor2 g18039(.a(new_n18232), .b(new_n18231), .O(new_n18233));
  inv1 g18040(.a(new_n18233), .O(new_n18234));
  nor2 g18041(.a(new_n17980), .b(new_n17855), .O(new_n18235));
  nor2 g18042(.a(new_n18235), .b(new_n18234), .O(new_n18236));
  inv1 g18043(.a(new_n18235), .O(new_n18237));
  nor2 g18044(.a(new_n18237), .b(new_n18233), .O(new_n18238));
  nor2 g18045(.a(new_n18238), .b(new_n18236), .O(new_n18239));
  nor2 g18046(.a(new_n17991), .b(new_n17987), .O(new_n18240));
  inv1 g18047(.a(new_n18240), .O(new_n18241));
  nor2 g18048(.a(new_n18241), .b(new_n18239), .O(new_n18242));
  inv1 g18049(.a(new_n18239), .O(new_n18243));
  nor2 g18050(.a(new_n18240), .b(new_n18243), .O(new_n18244));
  nor2 g18051(.a(new_n18244), .b(new_n18242), .O(new_n18245));
  inv1 g18052(.a(new_n18245), .O(\asquared[85] ));
  nor2 g18053(.a(new_n18231), .b(new_n18227), .O(new_n18247));
  nor2 g18054(.a(new_n18038), .b(new_n18032), .O(new_n18248));
  inv1 g18055(.a(new_n18248), .O(new_n18249));
  nor2 g18056(.a(new_n18101), .b(new_n18095), .O(new_n18250));
  inv1 g18057(.a(new_n18250), .O(new_n18251));
  nor2 g18058(.a(new_n18015), .b(new_n18009), .O(new_n18252));
  inv1 g18059(.a(new_n18252), .O(new_n18253));
  nor2 g18060(.a(new_n18253), .b(new_n18251), .O(new_n18254));
  nor2 g18061(.a(new_n18252), .b(new_n18250), .O(new_n18255));
  nor2 g18062(.a(new_n18255), .b(new_n18254), .O(new_n18256));
  nor2 g18063(.a(new_n18069), .b(new_n18053), .O(new_n18257));
  inv1 g18064(.a(new_n18257), .O(new_n18258));
  nor2 g18065(.a(new_n18258), .b(new_n18256), .O(new_n18259));
  inv1 g18066(.a(new_n18256), .O(new_n18260));
  nor2 g18067(.a(new_n18257), .b(new_n18260), .O(new_n18261));
  nor2 g18068(.a(new_n18261), .b(new_n18259), .O(new_n18262));
  nor2 g18069(.a(new_n18081), .b(new_n18075), .O(new_n18263));
  inv1 g18070(.a(new_n18263), .O(new_n18264));
  nor2 g18071(.a(new_n18264), .b(new_n18262), .O(new_n18265));
  inv1 g18072(.a(new_n18262), .O(new_n18266));
  nor2 g18073(.a(new_n18263), .b(new_n18266), .O(new_n18267));
  nor2 g18074(.a(new_n18267), .b(new_n18265), .O(new_n18268));
  inv1 g18075(.a(new_n18268), .O(new_n18269));
  nor2 g18076(.a(new_n18217), .b(new_n18213), .O(new_n18270));
  nor2 g18077(.a(new_n18270), .b(new_n18269), .O(new_n18271));
  inv1 g18078(.a(new_n18270), .O(new_n18272));
  nor2 g18079(.a(new_n18272), .b(new_n18268), .O(new_n18273));
  nor2 g18080(.a(new_n18273), .b(new_n18271), .O(new_n18274));
  nor2 g18081(.a(new_n18274), .b(new_n18249), .O(new_n18275));
  inv1 g18082(.a(new_n18274), .O(new_n18276));
  nor2 g18083(.a(new_n18276), .b(new_n18248), .O(new_n18277));
  nor2 g18084(.a(new_n18277), .b(new_n18275), .O(new_n18278));
  inv1 g18085(.a(new_n18278), .O(new_n18279));
  nor2 g18086(.a(new_n18221), .b(new_n18087), .O(new_n18280));
  nor2 g18087(.a(new_n18280), .b(new_n18279), .O(new_n18281));
  inv1 g18088(.a(new_n18280), .O(new_n18282));
  nor2 g18089(.a(new_n18282), .b(new_n18278), .O(new_n18283));
  nor2 g18090(.a(new_n18283), .b(new_n18281), .O(new_n18284));
  inv1 g18091(.a(new_n18284), .O(new_n18285));
  nor2 g18092(.a(new_n18042), .b(new_n18001), .O(new_n18286));
  nor2 g18093(.a(new_n18026), .b(new_n18023), .O(new_n18287));
  inv1 g18094(.a(new_n18287), .O(new_n18288));
  nor2 g18095(.a(new_n6274), .b(new_n4425), .O(new_n18289));
  inv1 g18096(.a(new_n18289), .O(new_n18290));
  nor2 g18097(.a(new_n5971), .b(new_n4682), .O(new_n18291));
  nor2 g18098(.a(new_n18291), .b(new_n18184), .O(new_n18292));
  nor2 g18099(.a(new_n5971), .b(new_n4954), .O(new_n18293));
  inv1 g18100(.a(new_n18293), .O(new_n18294));
  nor2 g18101(.a(new_n18294), .b(new_n17768), .O(new_n18295));
  nor2 g18102(.a(new_n18295), .b(new_n18292), .O(new_n18296));
  nor2 g18103(.a(new_n18296), .b(new_n18290), .O(new_n18297));
  inv1 g18104(.a(new_n18296), .O(new_n18298));
  nor2 g18105(.a(new_n18298), .b(new_n18289), .O(new_n18299));
  nor2 g18106(.a(new_n18299), .b(new_n18297), .O(new_n18300));
  nor2 g18107(.a(new_n8026), .b(new_n3231), .O(new_n18301));
  nor2 g18108(.a(new_n7537), .b(new_n3533), .O(new_n18302));
  nor2 g18109(.a(new_n18302), .b(new_n18301), .O(new_n18303));
  nor2 g18110(.a(new_n8026), .b(new_n3533), .O(new_n18304));
  inv1 g18111(.a(new_n18304), .O(new_n18305));
  nor2 g18112(.a(new_n18305), .b(new_n18145), .O(new_n18306));
  nor2 g18113(.a(new_n18306), .b(new_n18303), .O(new_n18307));
  nor2 g18114(.a(new_n18307), .b(new_n18062), .O(new_n18308));
  inv1 g18115(.a(new_n18307), .O(new_n18309));
  nor2 g18116(.a(new_n18309), .b(new_n18061), .O(new_n18310));
  nor2 g18117(.a(new_n18310), .b(new_n18308), .O(new_n18311));
  nor2 g18118(.a(new_n7294), .b(new_n3722), .O(new_n18312));
  inv1 g18119(.a(new_n18312), .O(new_n18313));
  nor2 g18120(.a(new_n9658), .b(new_n2433), .O(new_n18314));
  nor2 g18121(.a(new_n18314), .b(new_n17799), .O(new_n18315));
  inv1 g18122(.a(new_n18314), .O(new_n18316));
  nor2 g18123(.a(new_n18316), .b(new_n17800), .O(new_n18317));
  nor2 g18124(.a(new_n18317), .b(new_n18315), .O(new_n18318));
  inv1 g18125(.a(new_n18318), .O(new_n18319));
  nor2 g18126(.a(new_n18319), .b(new_n18313), .O(new_n18320));
  nor2 g18127(.a(new_n18318), .b(new_n18312), .O(new_n18321));
  nor2 g18128(.a(new_n18321), .b(new_n18320), .O(new_n18322));
  inv1 g18129(.a(new_n18322), .O(new_n18323));
  nor2 g18130(.a(new_n18323), .b(new_n18311), .O(new_n18324));
  inv1 g18131(.a(new_n18311), .O(new_n18325));
  nor2 g18132(.a(new_n18322), .b(new_n18325), .O(new_n18326));
  nor2 g18133(.a(new_n18326), .b(new_n18324), .O(new_n18327));
  nor2 g18134(.a(new_n18327), .b(new_n18300), .O(new_n18328));
  inv1 g18135(.a(new_n18300), .O(new_n18329));
  inv1 g18136(.a(new_n18327), .O(new_n18330));
  nor2 g18137(.a(new_n18330), .b(new_n18329), .O(new_n18331));
  nor2 g18138(.a(new_n18331), .b(new_n18328), .O(new_n18332));
  nor2 g18139(.a(new_n9156), .b(new_n2506), .O(new_n18333));
  inv1 g18140(.a(new_n18333), .O(new_n18334));
  nor2 g18141(.a(new_n8476), .b(new_n2826), .O(new_n18335));
  nor2 g18142(.a(new_n18335), .b(new_n17881), .O(new_n18336));
  inv1 g18143(.a(new_n18168), .O(new_n18337));
  nor2 g18144(.a(new_n8946), .b(new_n2826), .O(new_n18338));
  inv1 g18145(.a(new_n18338), .O(new_n18339));
  nor2 g18146(.a(new_n18339), .b(new_n18337), .O(new_n18340));
  nor2 g18147(.a(new_n18340), .b(new_n18336), .O(new_n18341));
  nor2 g18148(.a(new_n18341), .b(new_n18334), .O(new_n18342));
  inv1 g18149(.a(new_n18341), .O(new_n18343));
  nor2 g18150(.a(new_n18343), .b(new_n18333), .O(new_n18344));
  nor2 g18151(.a(new_n18344), .b(new_n18342), .O(new_n18345));
  inv1 g18152(.a(new_n18345), .O(new_n18346));
  nor2 g18153(.a(new_n6893), .b(new_n4093), .O(new_n18347));
  nor2 g18154(.a(new_n6570), .b(new_n4366), .O(new_n18348));
  nor2 g18155(.a(new_n18348), .b(new_n18347), .O(new_n18349));
  nor2 g18156(.a(new_n6893), .b(new_n4366), .O(new_n18350));
  inv1 g18157(.a(new_n18350), .O(new_n18351));
  nor2 g18158(.a(new_n18351), .b(new_n18167), .O(new_n18352));
  nor2 g18159(.a(new_n18352), .b(new_n18349), .O(new_n18353));
  nor2 g18160(.a(new_n18353), .b(new_n18122), .O(new_n18354));
  inv1 g18161(.a(new_n18353), .O(new_n18355));
  nor2 g18162(.a(new_n18355), .b(new_n18121), .O(new_n18356));
  nor2 g18163(.a(new_n18356), .b(new_n18354), .O(new_n18357));
  nor2 g18164(.a(new_n5393), .b(\a[42] ), .O(new_n18358));
  nor2 g18165(.a(new_n18358), .b(new_n18136), .O(new_n18359));
  inv1 g18166(.a(new_n18358), .O(new_n18360));
  nor2 g18167(.a(new_n18360), .b(new_n18135), .O(new_n18361));
  nor2 g18168(.a(new_n18361), .b(new_n18359), .O(new_n18362));
  nor2 g18169(.a(new_n18362), .b(new_n18357), .O(new_n18363));
  inv1 g18170(.a(new_n18357), .O(new_n18364));
  inv1 g18171(.a(new_n18362), .O(new_n18365));
  nor2 g18172(.a(new_n18365), .b(new_n18364), .O(new_n18366));
  nor2 g18173(.a(new_n18366), .b(new_n18363), .O(new_n18367));
  nor2 g18174(.a(new_n18367), .b(new_n18346), .O(new_n18368));
  inv1 g18175(.a(new_n18367), .O(new_n18369));
  nor2 g18176(.a(new_n18369), .b(new_n18345), .O(new_n18370));
  nor2 g18177(.a(new_n18370), .b(new_n18368), .O(new_n18371));
  inv1 g18178(.a(new_n18371), .O(new_n18372));
  nor2 g18179(.a(new_n18372), .b(new_n18332), .O(new_n18373));
  inv1 g18180(.a(new_n18332), .O(new_n18374));
  nor2 g18181(.a(new_n18371), .b(new_n18374), .O(new_n18375));
  nor2 g18182(.a(new_n18375), .b(new_n18373), .O(new_n18376));
  nor2 g18183(.a(new_n18376), .b(new_n18288), .O(new_n18377));
  inv1 g18184(.a(new_n18376), .O(new_n18378));
  nor2 g18185(.a(new_n18378), .b(new_n18287), .O(new_n18379));
  nor2 g18186(.a(new_n18379), .b(new_n18377), .O(new_n18380));
  inv1 g18187(.a(new_n18380), .O(new_n18381));
  nor2 g18188(.a(new_n18127), .b(new_n18119), .O(new_n18382));
  nor2 g18189(.a(new_n18140), .b(new_n18133), .O(new_n18383));
  nor2 g18190(.a(new_n18383), .b(new_n18382), .O(new_n18384));
  inv1 g18191(.a(new_n18382), .O(new_n18385));
  inv1 g18192(.a(new_n18383), .O(new_n18386));
  nor2 g18193(.a(new_n18386), .b(new_n18385), .O(new_n18387));
  nor2 g18194(.a(new_n18387), .b(new_n18384), .O(new_n18388));
  nor2 g18195(.a(new_n18154), .b(new_n18147), .O(new_n18389));
  nor2 g18196(.a(new_n18389), .b(new_n18388), .O(new_n18390));
  inv1 g18197(.a(new_n18388), .O(new_n18391));
  inv1 g18198(.a(new_n18389), .O(new_n18392));
  nor2 g18199(.a(new_n18392), .b(new_n18391), .O(new_n18393));
  nor2 g18200(.a(new_n18393), .b(new_n18390), .O(new_n18394));
  inv1 g18201(.a(new_n18394), .O(new_n18395));
  nor2 g18202(.a(new_n18210), .b(new_n18203), .O(new_n18396));
  inv1 g18203(.a(new_n18396), .O(new_n18397));
  nor2 g18204(.a(new_n18163), .b(new_n18156), .O(new_n18398));
  inv1 g18205(.a(new_n18398), .O(new_n18399));
  nor2 g18206(.a(new_n18399), .b(new_n18397), .O(new_n18400));
  nor2 g18207(.a(new_n18398), .b(new_n18396), .O(new_n18401));
  nor2 g18208(.a(new_n18401), .b(new_n18400), .O(new_n18402));
  inv1 g18209(.a(new_n18402), .O(new_n18403));
  nor2 g18210(.a(new_n18403), .b(new_n18395), .O(new_n18404));
  nor2 g18211(.a(new_n18402), .b(new_n18394), .O(new_n18405));
  nor2 g18212(.a(new_n18405), .b(new_n18404), .O(new_n18406));
  inv1 g18213(.a(new_n18406), .O(new_n18407));
  nor2 g18214(.a(new_n18112), .b(new_n18109), .O(new_n18408));
  nor2 g18215(.a(new_n10895), .b(new_n1736), .O(new_n18409));
  inv1 g18216(.a(new_n18409), .O(new_n18410));
  nor2 g18217(.a(new_n18190), .b(new_n18182), .O(new_n18411));
  inv1 g18218(.a(new_n18411), .O(new_n18412));
  nor2 g18219(.a(new_n18412), .b(new_n18410), .O(new_n18413));
  nor2 g18220(.a(new_n18411), .b(new_n18409), .O(new_n18414));
  nor2 g18221(.a(new_n18414), .b(new_n18413), .O(new_n18415));
  nor2 g18222(.a(new_n18201), .b(new_n18195), .O(new_n18416));
  nor2 g18223(.a(new_n18416), .b(new_n18415), .O(new_n18417));
  inv1 g18224(.a(new_n18415), .O(new_n18418));
  inv1 g18225(.a(new_n18416), .O(new_n18419));
  nor2 g18226(.a(new_n18419), .b(new_n18418), .O(new_n18420));
  nor2 g18227(.a(new_n18420), .b(new_n18417), .O(new_n18421));
  inv1 g18228(.a(new_n18421), .O(new_n18422));
  nor2 g18229(.a(new_n18067), .b(new_n18060), .O(new_n18423));
  nor2 g18230(.a(new_n18176), .b(new_n18169), .O(new_n18424));
  nor2 g18231(.a(new_n18424), .b(new_n18423), .O(new_n18425));
  inv1 g18232(.a(new_n18423), .O(new_n18426));
  inv1 g18233(.a(new_n18424), .O(new_n18427));
  nor2 g18234(.a(new_n18427), .b(new_n18426), .O(new_n18428));
  nor2 g18235(.a(new_n18428), .b(new_n18425), .O(new_n18429));
  inv1 g18236(.a(new_n18429), .O(new_n18430));
  nor2 g18237(.a(new_n10320), .b(new_n2121), .O(new_n18431));
  nor2 g18238(.a(new_n9873), .b(new_n2184), .O(new_n18432));
  nor2 g18239(.a(new_n18432), .b(new_n18431), .O(new_n18433));
  nor2 g18240(.a(new_n18057), .b(new_n10325), .O(new_n18434));
  nor2 g18241(.a(new_n18434), .b(new_n18433), .O(new_n18435));
  nor2 g18242(.a(new_n18435), .b(new_n18149), .O(new_n18436));
  inv1 g18243(.a(new_n18435), .O(new_n18437));
  nor2 g18244(.a(new_n18437), .b(new_n18148), .O(new_n18438));
  nor2 g18245(.a(new_n18438), .b(new_n18436), .O(new_n18439));
  nor2 g18246(.a(new_n18439), .b(new_n18430), .O(new_n18440));
  inv1 g18247(.a(new_n18439), .O(new_n18441));
  nor2 g18248(.a(new_n18441), .b(new_n18429), .O(new_n18442));
  nor2 g18249(.a(new_n18442), .b(new_n18440), .O(new_n18443));
  inv1 g18250(.a(new_n18443), .O(new_n18444));
  nor2 g18251(.a(new_n18444), .b(new_n18422), .O(new_n18445));
  nor2 g18252(.a(new_n18443), .b(new_n18421), .O(new_n18446));
  nor2 g18253(.a(new_n18446), .b(new_n18445), .O(new_n18447));
  inv1 g18254(.a(new_n18447), .O(new_n18448));
  nor2 g18255(.a(new_n18448), .b(new_n18408), .O(new_n18449));
  inv1 g18256(.a(new_n18408), .O(new_n18450));
  nor2 g18257(.a(new_n18447), .b(new_n18450), .O(new_n18451));
  nor2 g18258(.a(new_n18451), .b(new_n18449), .O(new_n18452));
  inv1 g18259(.a(new_n18452), .O(new_n18453));
  nor2 g18260(.a(new_n18453), .b(new_n18407), .O(new_n18454));
  nor2 g18261(.a(new_n18452), .b(new_n18406), .O(new_n18455));
  nor2 g18262(.a(new_n18455), .b(new_n18454), .O(new_n18456));
  inv1 g18263(.a(new_n18456), .O(new_n18457));
  nor2 g18264(.a(new_n18457), .b(new_n18381), .O(new_n18458));
  nor2 g18265(.a(new_n18456), .b(new_n18380), .O(new_n18459));
  nor2 g18266(.a(new_n18459), .b(new_n18458), .O(new_n18460));
  inv1 g18267(.a(new_n18460), .O(new_n18461));
  nor2 g18268(.a(new_n18461), .b(new_n18286), .O(new_n18462));
  inv1 g18269(.a(new_n18286), .O(new_n18463));
  nor2 g18270(.a(new_n18460), .b(new_n18463), .O(new_n18464));
  nor2 g18271(.a(new_n18464), .b(new_n18462), .O(new_n18465));
  inv1 g18272(.a(new_n18465), .O(new_n18466));
  nor2 g18273(.a(new_n18466), .b(new_n18285), .O(new_n18467));
  nor2 g18274(.a(new_n18465), .b(new_n18284), .O(new_n18468));
  nor2 g18275(.a(new_n18468), .b(new_n18467), .O(new_n18469));
  inv1 g18276(.a(new_n18469), .O(new_n18470));
  nor2 g18277(.a(new_n18470), .b(new_n18247), .O(new_n18471));
  inv1 g18278(.a(new_n18247), .O(new_n18472));
  nor2 g18279(.a(new_n18469), .b(new_n18472), .O(new_n18473));
  nor2 g18280(.a(new_n18473), .b(new_n18471), .O(new_n18474));
  inv1 g18281(.a(new_n18474), .O(new_n18475));
  nor2 g18282(.a(new_n18240), .b(new_n18236), .O(new_n18476));
  nor2 g18283(.a(new_n18476), .b(new_n18238), .O(new_n18477));
  nor2 g18284(.a(new_n18477), .b(new_n18475), .O(new_n18478));
  inv1 g18285(.a(new_n18477), .O(new_n18479));
  nor2 g18286(.a(new_n18479), .b(new_n18474), .O(new_n18480));
  nor2 g18287(.a(new_n18480), .b(new_n18478), .O(new_n18481));
  inv1 g18288(.a(new_n18481), .O(\asquared[86] ));
  nor2 g18289(.a(new_n18467), .b(new_n18462), .O(new_n18483));
  inv1 g18290(.a(new_n18483), .O(new_n18484));
  nor2 g18291(.a(new_n18458), .b(new_n18454), .O(new_n18485));
  inv1 g18292(.a(new_n18485), .O(new_n18486));
  nor2 g18293(.a(new_n18271), .b(new_n18267), .O(new_n18487));
  inv1 g18294(.a(new_n18487), .O(new_n18488));
  nor2 g18295(.a(new_n18488), .b(new_n18486), .O(new_n18489));
  nor2 g18296(.a(new_n18487), .b(new_n18485), .O(new_n18490));
  nor2 g18297(.a(new_n18490), .b(new_n18489), .O(new_n18491));
  inv1 g18298(.a(new_n18491), .O(new_n18492));
  nor2 g18299(.a(new_n18449), .b(new_n18445), .O(new_n18493));
  nor2 g18300(.a(new_n18420), .b(new_n18413), .O(new_n18494));
  inv1 g18301(.a(new_n18494), .O(new_n18495));
  nor2 g18302(.a(new_n10895), .b(new_n1903), .O(new_n18496));
  nor2 g18303(.a(new_n11186), .b(new_n1736), .O(new_n18497));
  nor2 g18304(.a(new_n18497), .b(new_n18496), .O(new_n18498));
  nor2 g18305(.a(new_n11186), .b(new_n1903), .O(new_n18499));
  inv1 g18306(.a(new_n18499), .O(new_n18500));
  nor2 g18307(.a(new_n18500), .b(new_n18410), .O(new_n18501));
  nor2 g18308(.a(new_n18501), .b(new_n18498), .O(new_n18502));
  inv1 g18309(.a(new_n18502), .O(new_n18503));
  nor2 g18310(.a(new_n18361), .b(new_n5393), .O(new_n18504));
  inv1 g18311(.a(new_n18504), .O(new_n18505));
  nor2 g18312(.a(new_n18505), .b(new_n18503), .O(new_n18506));
  nor2 g18313(.a(new_n18504), .b(new_n18502), .O(new_n18507));
  nor2 g18314(.a(new_n18507), .b(new_n18506), .O(new_n18508));
  nor2 g18315(.a(new_n18508), .b(new_n18495), .O(new_n18509));
  inv1 g18316(.a(new_n18508), .O(new_n18510));
  nor2 g18317(.a(new_n18510), .b(new_n18494), .O(new_n18511));
  nor2 g18318(.a(new_n18511), .b(new_n18509), .O(new_n18512));
  nor2 g18319(.a(new_n18393), .b(new_n18387), .O(new_n18513));
  inv1 g18320(.a(new_n18513), .O(new_n18514));
  nor2 g18321(.a(new_n18514), .b(new_n18512), .O(new_n18515));
  inv1 g18322(.a(new_n18512), .O(new_n18516));
  nor2 g18323(.a(new_n18513), .b(new_n18516), .O(new_n18517));
  nor2 g18324(.a(new_n18517), .b(new_n18515), .O(new_n18518));
  inv1 g18325(.a(new_n18518), .O(new_n18519));
  nor2 g18326(.a(new_n18519), .b(new_n18493), .O(new_n18520));
  inv1 g18327(.a(new_n18493), .O(new_n18521));
  nor2 g18328(.a(new_n18518), .b(new_n18521), .O(new_n18522));
  nor2 g18329(.a(new_n18522), .b(new_n18520), .O(new_n18523));
  inv1 g18330(.a(new_n18523), .O(new_n18524));
  nor2 g18331(.a(new_n18379), .b(new_n18373), .O(new_n18525));
  nor2 g18332(.a(new_n18525), .b(new_n18524), .O(new_n18526));
  inv1 g18333(.a(new_n18525), .O(new_n18527));
  nor2 g18334(.a(new_n18527), .b(new_n18523), .O(new_n18528));
  nor2 g18335(.a(new_n18528), .b(new_n18526), .O(new_n18529));
  inv1 g18336(.a(new_n18529), .O(new_n18530));
  nor2 g18337(.a(new_n18530), .b(new_n18492), .O(new_n18531));
  nor2 g18338(.a(new_n18529), .b(new_n18491), .O(new_n18532));
  nor2 g18339(.a(new_n18532), .b(new_n18531), .O(new_n18533));
  inv1 g18340(.a(new_n18533), .O(new_n18534));
  nor2 g18341(.a(new_n18281), .b(new_n18277), .O(new_n18535));
  nor2 g18342(.a(new_n18440), .b(new_n18428), .O(new_n18536));
  inv1 g18343(.a(new_n18536), .O(new_n18537));
  nor2 g18344(.a(new_n18331), .b(new_n18326), .O(new_n18538));
  nor2 g18345(.a(new_n18538), .b(new_n18537), .O(new_n18539));
  inv1 g18346(.a(new_n18538), .O(new_n18540));
  nor2 g18347(.a(new_n18540), .b(new_n18536), .O(new_n18541));
  nor2 g18348(.a(new_n18541), .b(new_n18539), .O(new_n18542));
  nor2 g18349(.a(new_n18370), .b(new_n18363), .O(new_n18543));
  inv1 g18350(.a(new_n18543), .O(new_n18544));
  nor2 g18351(.a(new_n18544), .b(new_n18542), .O(new_n18545));
  inv1 g18352(.a(new_n18542), .O(new_n18546));
  nor2 g18353(.a(new_n18543), .b(new_n18546), .O(new_n18547));
  nor2 g18354(.a(new_n18547), .b(new_n18545), .O(new_n18548));
  inv1 g18355(.a(new_n18548), .O(new_n18549));
  nor2 g18356(.a(new_n18261), .b(new_n18255), .O(new_n18550));
  nor2 g18357(.a(new_n18299), .b(new_n18292), .O(new_n18551));
  nor2 g18358(.a(new_n18344), .b(new_n18336), .O(new_n18552));
  nor2 g18359(.a(new_n18552), .b(new_n18551), .O(new_n18553));
  inv1 g18360(.a(new_n18551), .O(new_n18554));
  inv1 g18361(.a(new_n18552), .O(new_n18555));
  nor2 g18362(.a(new_n18555), .b(new_n18554), .O(new_n18556));
  nor2 g18363(.a(new_n18556), .b(new_n18553), .O(new_n18557));
  nor2 g18364(.a(new_n18356), .b(new_n18349), .O(new_n18558));
  nor2 g18365(.a(new_n18558), .b(new_n18557), .O(new_n18559));
  inv1 g18366(.a(new_n18557), .O(new_n18560));
  inv1 g18367(.a(new_n18558), .O(new_n18561));
  nor2 g18368(.a(new_n18561), .b(new_n18560), .O(new_n18562));
  nor2 g18369(.a(new_n18562), .b(new_n18559), .O(new_n18563));
  inv1 g18370(.a(new_n18563), .O(new_n18564));
  nor2 g18371(.a(new_n18320), .b(new_n18317), .O(new_n18565));
  inv1 g18372(.a(new_n18565), .O(new_n18566));
  nor2 g18373(.a(new_n18310), .b(new_n18303), .O(new_n18567));
  nor2 g18374(.a(new_n18438), .b(new_n18433), .O(new_n18568));
  nor2 g18375(.a(new_n18568), .b(new_n18567), .O(new_n18569));
  inv1 g18376(.a(new_n18567), .O(new_n18570));
  inv1 g18377(.a(new_n18568), .O(new_n18571));
  nor2 g18378(.a(new_n18571), .b(new_n18570), .O(new_n18572));
  nor2 g18379(.a(new_n18572), .b(new_n18569), .O(new_n18573));
  nor2 g18380(.a(new_n18573), .b(new_n18566), .O(new_n18574));
  inv1 g18381(.a(new_n18573), .O(new_n18575));
  nor2 g18382(.a(new_n18575), .b(new_n18565), .O(new_n18576));
  nor2 g18383(.a(new_n18576), .b(new_n18574), .O(new_n18577));
  inv1 g18384(.a(new_n18577), .O(new_n18578));
  nor2 g18385(.a(new_n18578), .b(new_n18564), .O(new_n18579));
  nor2 g18386(.a(new_n18577), .b(new_n18563), .O(new_n18580));
  nor2 g18387(.a(new_n18580), .b(new_n18579), .O(new_n18581));
  inv1 g18388(.a(new_n18581), .O(new_n18582));
  nor2 g18389(.a(new_n18582), .b(new_n18550), .O(new_n18583));
  inv1 g18390(.a(new_n18550), .O(new_n18584));
  nor2 g18391(.a(new_n18581), .b(new_n18584), .O(new_n18585));
  nor2 g18392(.a(new_n18585), .b(new_n18583), .O(new_n18586));
  inv1 g18393(.a(new_n18586), .O(new_n18587));
  nor2 g18394(.a(new_n18587), .b(new_n18549), .O(new_n18588));
  nor2 g18395(.a(new_n18586), .b(new_n18548), .O(new_n18589));
  nor2 g18396(.a(new_n18589), .b(new_n18588), .O(new_n18590));
  inv1 g18397(.a(new_n18590), .O(new_n18591));
  nor2 g18398(.a(new_n18404), .b(new_n18401), .O(new_n18592));
  nor2 g18399(.a(new_n9156), .b(new_n2660), .O(new_n18593));
  inv1 g18400(.a(new_n18593), .O(new_n18594));
  nor2 g18401(.a(new_n6274), .b(new_n4682), .O(new_n18595));
  nor2 g18402(.a(new_n6570), .b(new_n4425), .O(new_n18596));
  nor2 g18403(.a(new_n18596), .b(new_n18595), .O(new_n18597));
  nor2 g18404(.a(new_n6570), .b(new_n4682), .O(new_n18598));
  inv1 g18405(.a(new_n18598), .O(new_n18599));
  nor2 g18406(.a(new_n18599), .b(new_n18290), .O(new_n18600));
  nor2 g18407(.a(new_n18600), .b(new_n18597), .O(new_n18601));
  nor2 g18408(.a(new_n18601), .b(new_n18594), .O(new_n18602));
  inv1 g18409(.a(new_n18601), .O(new_n18603));
  nor2 g18410(.a(new_n18603), .b(new_n18593), .O(new_n18604));
  nor2 g18411(.a(new_n18604), .b(new_n18602), .O(new_n18605));
  nor2 g18412(.a(new_n10468), .b(new_n2121), .O(new_n18606));
  nor2 g18413(.a(new_n9873), .b(new_n2433), .O(new_n18607));
  nor2 g18414(.a(new_n18607), .b(new_n10324), .O(new_n18608));
  inv1 g18415(.a(new_n18432), .O(new_n18609));
  nor2 g18416(.a(new_n10320), .b(new_n2433), .O(new_n18610));
  inv1 g18417(.a(new_n18610), .O(new_n18611));
  nor2 g18418(.a(new_n18611), .b(new_n18609), .O(new_n18612));
  nor2 g18419(.a(new_n18612), .b(new_n18608), .O(new_n18613));
  inv1 g18420(.a(new_n18613), .O(new_n18614));
  nor2 g18421(.a(new_n18614), .b(new_n18606), .O(new_n18615));
  inv1 g18422(.a(new_n18606), .O(new_n18616));
  nor2 g18423(.a(new_n18613), .b(new_n18616), .O(new_n18617));
  nor2 g18424(.a(new_n18617), .b(new_n18615), .O(new_n18618));
  nor2 g18425(.a(new_n8476), .b(new_n3057), .O(new_n18619));
  nor2 g18426(.a(new_n5796), .b(new_n5178), .O(new_n18620));
  nor2 g18427(.a(new_n18620), .b(new_n18619), .O(new_n18621));
  inv1 g18428(.a(new_n18619), .O(new_n18622));
  inv1 g18429(.a(new_n18620), .O(new_n18623));
  nor2 g18430(.a(new_n18623), .b(new_n18622), .O(new_n18624));
  nor2 g18431(.a(new_n18624), .b(new_n18621), .O(new_n18625));
  nor2 g18432(.a(new_n18625), .b(new_n18294), .O(new_n18626));
  inv1 g18433(.a(new_n18625), .O(new_n18627));
  nor2 g18434(.a(new_n18627), .b(new_n18293), .O(new_n18628));
  nor2 g18435(.a(new_n18628), .b(new_n18626), .O(new_n18629));
  nor2 g18436(.a(new_n18629), .b(new_n18618), .O(new_n18630));
  inv1 g18437(.a(new_n18618), .O(new_n18631));
  inv1 g18438(.a(new_n18629), .O(new_n18632));
  nor2 g18439(.a(new_n18632), .b(new_n18631), .O(new_n18633));
  nor2 g18440(.a(new_n18633), .b(new_n18630), .O(new_n18634));
  inv1 g18441(.a(new_n18634), .O(new_n18635));
  nor2 g18442(.a(new_n18635), .b(new_n18605), .O(new_n18636));
  inv1 g18443(.a(new_n18605), .O(new_n18637));
  nor2 g18444(.a(new_n18634), .b(new_n18637), .O(new_n18638));
  nor2 g18445(.a(new_n18638), .b(new_n18636), .O(new_n18639));
  nor2 g18446(.a(new_n9658), .b(new_n2506), .O(new_n18640));
  nor2 g18447(.a(new_n18640), .b(new_n18338), .O(new_n18641));
  nor2 g18448(.a(new_n9658), .b(new_n2826), .O(new_n18642));
  inv1 g18449(.a(new_n18642), .O(new_n18643));
  nor2 g18450(.a(new_n18643), .b(new_n18196), .O(new_n18644));
  nor2 g18451(.a(new_n18644), .b(new_n18641), .O(new_n18645));
  nor2 g18452(.a(new_n18645), .b(new_n18351), .O(new_n18646));
  inv1 g18453(.a(new_n18645), .O(new_n18647));
  nor2 g18454(.a(new_n18647), .b(new_n18350), .O(new_n18648));
  nor2 g18455(.a(new_n18648), .b(new_n18646), .O(new_n18649));
  inv1 g18456(.a(new_n18649), .O(new_n18650));
  nor2 g18457(.a(new_n11596), .b(new_n1647), .O(new_n18651));
  nor2 g18458(.a(new_n7294), .b(new_n3870), .O(new_n18652));
  nor2 g18459(.a(new_n6958), .b(new_n4093), .O(new_n18653));
  nor2 g18460(.a(new_n18653), .b(new_n18652), .O(new_n18654));
  nor2 g18461(.a(new_n7294), .b(new_n4093), .O(new_n18655));
  inv1 g18462(.a(new_n18655), .O(new_n18656));
  nor2 g18463(.a(new_n18656), .b(new_n18122), .O(new_n18657));
  nor2 g18464(.a(new_n18657), .b(new_n18654), .O(new_n18658));
  inv1 g18465(.a(new_n18658), .O(new_n18659));
  nor2 g18466(.a(new_n18659), .b(new_n18651), .O(new_n18660));
  inv1 g18467(.a(new_n18651), .O(new_n18661));
  nor2 g18468(.a(new_n18658), .b(new_n18661), .O(new_n18662));
  nor2 g18469(.a(new_n18662), .b(new_n18660), .O(new_n18663));
  nor2 g18470(.a(new_n8170), .b(new_n3231), .O(new_n18664));
  inv1 g18471(.a(new_n18664), .O(new_n18665));
  nor2 g18472(.a(new_n7537), .b(new_n3722), .O(new_n18666));
  nor2 g18473(.a(new_n18666), .b(new_n18304), .O(new_n18667));
  inv1 g18474(.a(new_n18302), .O(new_n18668));
  nor2 g18475(.a(new_n8026), .b(new_n3722), .O(new_n18669));
  inv1 g18476(.a(new_n18669), .O(new_n18670));
  nor2 g18477(.a(new_n18670), .b(new_n18668), .O(new_n18671));
  nor2 g18478(.a(new_n18671), .b(new_n18667), .O(new_n18672));
  nor2 g18479(.a(new_n18672), .b(new_n18665), .O(new_n18673));
  inv1 g18480(.a(new_n18672), .O(new_n18674));
  nor2 g18481(.a(new_n18674), .b(new_n18664), .O(new_n18675));
  nor2 g18482(.a(new_n18675), .b(new_n18673), .O(new_n18676));
  nor2 g18483(.a(new_n18676), .b(new_n18663), .O(new_n18677));
  inv1 g18484(.a(new_n18663), .O(new_n18678));
  inv1 g18485(.a(new_n18676), .O(new_n18679));
  nor2 g18486(.a(new_n18679), .b(new_n18678), .O(new_n18680));
  nor2 g18487(.a(new_n18680), .b(new_n18677), .O(new_n18681));
  nor2 g18488(.a(new_n18681), .b(new_n18650), .O(new_n18682));
  inv1 g18489(.a(new_n18681), .O(new_n18683));
  nor2 g18490(.a(new_n18683), .b(new_n18649), .O(new_n18684));
  nor2 g18491(.a(new_n18684), .b(new_n18682), .O(new_n18685));
  nor2 g18492(.a(new_n18685), .b(new_n18639), .O(new_n18686));
  inv1 g18493(.a(new_n18639), .O(new_n18687));
  inv1 g18494(.a(new_n18685), .O(new_n18688));
  nor2 g18495(.a(new_n18688), .b(new_n18687), .O(new_n18689));
  nor2 g18496(.a(new_n18689), .b(new_n18686), .O(new_n18690));
  inv1 g18497(.a(new_n18690), .O(new_n18691));
  nor2 g18498(.a(new_n18691), .b(new_n18592), .O(new_n18692));
  inv1 g18499(.a(new_n18592), .O(new_n18693));
  nor2 g18500(.a(new_n18690), .b(new_n18693), .O(new_n18694));
  nor2 g18501(.a(new_n18694), .b(new_n18692), .O(new_n18695));
  inv1 g18502(.a(new_n18695), .O(new_n18696));
  nor2 g18503(.a(new_n18696), .b(new_n18591), .O(new_n18697));
  nor2 g18504(.a(new_n18695), .b(new_n18590), .O(new_n18698));
  nor2 g18505(.a(new_n18698), .b(new_n18697), .O(new_n18699));
  inv1 g18506(.a(new_n18699), .O(new_n18700));
  nor2 g18507(.a(new_n18700), .b(new_n18535), .O(new_n18701));
  inv1 g18508(.a(new_n18535), .O(new_n18702));
  nor2 g18509(.a(new_n18699), .b(new_n18702), .O(new_n18703));
  nor2 g18510(.a(new_n18703), .b(new_n18701), .O(new_n18704));
  inv1 g18511(.a(new_n18704), .O(new_n18705));
  nor2 g18512(.a(new_n18705), .b(new_n18534), .O(new_n18706));
  nor2 g18513(.a(new_n18704), .b(new_n18533), .O(new_n18707));
  nor2 g18514(.a(new_n18707), .b(new_n18706), .O(new_n18708));
  nor2 g18515(.a(new_n18708), .b(new_n18484), .O(new_n18709));
  inv1 g18516(.a(new_n18708), .O(new_n18710));
  nor2 g18517(.a(new_n18710), .b(new_n18483), .O(new_n18711));
  nor2 g18518(.a(new_n18711), .b(new_n18709), .O(new_n18712));
  nor2 g18519(.a(new_n18478), .b(new_n18473), .O(new_n18713));
  inv1 g18520(.a(new_n18713), .O(new_n18714));
  nor2 g18521(.a(new_n18714), .b(new_n18712), .O(new_n18715));
  inv1 g18522(.a(new_n18712), .O(new_n18716));
  nor2 g18523(.a(new_n18713), .b(new_n18716), .O(new_n18717));
  nor2 g18524(.a(new_n18717), .b(new_n18715), .O(new_n18718));
  inv1 g18525(.a(new_n18718), .O(\asquared[87] ));
  nor2 g18526(.a(new_n18706), .b(new_n18701), .O(new_n18720));
  inv1 g18527(.a(new_n18720), .O(new_n18721));
  nor2 g18528(.a(new_n18692), .b(new_n18689), .O(new_n18722));
  nor2 g18529(.a(new_n18562), .b(new_n18556), .O(new_n18723));
  inv1 g18530(.a(new_n18723), .O(new_n18724));
  nor2 g18531(.a(new_n18684), .b(new_n18677), .O(new_n18725));
  inv1 g18532(.a(new_n18725), .O(new_n18726));
  nor2 g18533(.a(new_n18726), .b(new_n18724), .O(new_n18727));
  nor2 g18534(.a(new_n18725), .b(new_n18723), .O(new_n18728));
  nor2 g18535(.a(new_n18728), .b(new_n18727), .O(new_n18729));
  nor2 g18536(.a(new_n18636), .b(new_n18630), .O(new_n18730));
  inv1 g18537(.a(new_n18730), .O(new_n18731));
  nor2 g18538(.a(new_n18731), .b(new_n18729), .O(new_n18732));
  inv1 g18539(.a(new_n18729), .O(new_n18733));
  nor2 g18540(.a(new_n18730), .b(new_n18733), .O(new_n18734));
  nor2 g18541(.a(new_n18734), .b(new_n18732), .O(new_n18735));
  inv1 g18542(.a(new_n18735), .O(new_n18736));
  nor2 g18543(.a(new_n18736), .b(new_n18722), .O(new_n18737));
  inv1 g18544(.a(new_n18722), .O(new_n18738));
  nor2 g18545(.a(new_n18735), .b(new_n18738), .O(new_n18739));
  nor2 g18546(.a(new_n18739), .b(new_n18737), .O(new_n18740));
  nor2 g18547(.a(new_n18526), .b(new_n18520), .O(new_n18741));
  inv1 g18548(.a(new_n18741), .O(new_n18742));
  nor2 g18549(.a(new_n18742), .b(new_n18740), .O(new_n18743));
  inv1 g18550(.a(new_n18740), .O(new_n18744));
  nor2 g18551(.a(new_n18741), .b(new_n18744), .O(new_n18745));
  nor2 g18552(.a(new_n18745), .b(new_n18743), .O(new_n18746));
  nor2 g18553(.a(new_n18531), .b(new_n18490), .O(new_n18747));
  inv1 g18554(.a(new_n18747), .O(new_n18748));
  nor2 g18555(.a(new_n18748), .b(new_n18746), .O(new_n18749));
  inv1 g18556(.a(new_n18746), .O(new_n18750));
  nor2 g18557(.a(new_n18747), .b(new_n18750), .O(new_n18751));
  nor2 g18558(.a(new_n18751), .b(new_n18749), .O(new_n18752));
  nor2 g18559(.a(new_n18697), .b(new_n18588), .O(new_n18753));
  nor2 g18560(.a(new_n18576), .b(new_n18572), .O(new_n18754));
  inv1 g18561(.a(new_n18754), .O(new_n18755));
  nor2 g18562(.a(new_n9156), .b(new_n2826), .O(new_n18756));
  nor2 g18563(.a(new_n8476), .b(new_n3231), .O(new_n18757));
  nor2 g18564(.a(new_n18757), .b(new_n18756), .O(new_n18758));
  inv1 g18565(.a(new_n18335), .O(new_n18759));
  nor2 g18566(.a(new_n9156), .b(new_n3231), .O(new_n18760));
  inv1 g18567(.a(new_n18760), .O(new_n18761));
  nor2 g18568(.a(new_n18761), .b(new_n18759), .O(new_n18762));
  nor2 g18569(.a(new_n18762), .b(new_n18758), .O(new_n18763));
  nor2 g18570(.a(new_n18763), .b(new_n18599), .O(new_n18764));
  inv1 g18571(.a(new_n18763), .O(new_n18765));
  nor2 g18572(.a(new_n18765), .b(new_n18598), .O(new_n18766));
  nor2 g18573(.a(new_n18766), .b(new_n18764), .O(new_n18767));
  nor2 g18574(.a(new_n5796), .b(\a[43] ), .O(new_n18768));
  nor2 g18575(.a(new_n18768), .b(new_n18500), .O(new_n18769));
  inv1 g18576(.a(new_n18768), .O(new_n18770));
  nor2 g18577(.a(new_n18770), .b(new_n18499), .O(new_n18771));
  nor2 g18578(.a(new_n18771), .b(new_n18769), .O(new_n18772));
  nor2 g18579(.a(new_n18772), .b(new_n18767), .O(new_n18773));
  inv1 g18580(.a(new_n18767), .O(new_n18774));
  inv1 g18581(.a(new_n18772), .O(new_n18775));
  nor2 g18582(.a(new_n18775), .b(new_n18774), .O(new_n18776));
  nor2 g18583(.a(new_n18776), .b(new_n18773), .O(new_n18777));
  nor2 g18584(.a(new_n18777), .b(new_n18755), .O(new_n18778));
  inv1 g18585(.a(new_n18777), .O(new_n18779));
  nor2 g18586(.a(new_n18779), .b(new_n18754), .O(new_n18780));
  nor2 g18587(.a(new_n18780), .b(new_n18778), .O(new_n18781));
  nor2 g18588(.a(new_n8946), .b(new_n3057), .O(new_n18782));
  inv1 g18589(.a(new_n18782), .O(new_n18783));
  nor2 g18590(.a(new_n5971), .b(new_n5178), .O(new_n18784));
  nor2 g18591(.a(new_n6274), .b(new_n4954), .O(new_n18785));
  nor2 g18592(.a(new_n18785), .b(new_n18784), .O(new_n18786));
  nor2 g18593(.a(new_n6274), .b(new_n5178), .O(new_n18787));
  inv1 g18594(.a(new_n18787), .O(new_n18788));
  nor2 g18595(.a(new_n18788), .b(new_n18294), .O(new_n18789));
  nor2 g18596(.a(new_n18789), .b(new_n18786), .O(new_n18790));
  nor2 g18597(.a(new_n18790), .b(new_n18783), .O(new_n18791));
  inv1 g18598(.a(new_n18790), .O(new_n18792));
  nor2 g18599(.a(new_n18792), .b(new_n18782), .O(new_n18793));
  nor2 g18600(.a(new_n18793), .b(new_n18791), .O(new_n18794));
  inv1 g18601(.a(new_n18794), .O(new_n18795));
  nor2 g18602(.a(new_n11596), .b(new_n1736), .O(new_n18796));
  nor2 g18603(.a(new_n10895), .b(new_n2121), .O(new_n18797));
  nor2 g18604(.a(new_n10468), .b(new_n2184), .O(new_n18798));
  nor2 g18605(.a(new_n18798), .b(new_n18797), .O(new_n18799));
  nor2 g18606(.a(new_n10895), .b(new_n2184), .O(new_n18800));
  inv1 g18607(.a(new_n18800), .O(new_n18801));
  nor2 g18608(.a(new_n18801), .b(new_n18616), .O(new_n18802));
  nor2 g18609(.a(new_n18802), .b(new_n18799), .O(new_n18803));
  inv1 g18610(.a(new_n18803), .O(new_n18804));
  nor2 g18611(.a(new_n18804), .b(new_n18796), .O(new_n18805));
  inv1 g18612(.a(new_n18796), .O(new_n18806));
  nor2 g18613(.a(new_n18803), .b(new_n18806), .O(new_n18807));
  nor2 g18614(.a(new_n18807), .b(new_n18805), .O(new_n18808));
  nor2 g18615(.a(new_n6958), .b(new_n4366), .O(new_n18809));
  nor2 g18616(.a(new_n6893), .b(new_n4425), .O(new_n18810));
  nor2 g18617(.a(new_n18810), .b(new_n18809), .O(new_n18811));
  nor2 g18618(.a(new_n6958), .b(new_n4425), .O(new_n18812));
  inv1 g18619(.a(new_n18812), .O(new_n18813));
  nor2 g18620(.a(new_n18813), .b(new_n18351), .O(new_n18814));
  nor2 g18621(.a(new_n18814), .b(new_n18811), .O(new_n18815));
  nor2 g18622(.a(new_n18815), .b(new_n18656), .O(new_n18816));
  inv1 g18623(.a(new_n18815), .O(new_n18817));
  nor2 g18624(.a(new_n18817), .b(new_n18655), .O(new_n18818));
  nor2 g18625(.a(new_n18818), .b(new_n18816), .O(new_n18819));
  nor2 g18626(.a(new_n18819), .b(new_n18808), .O(new_n18820));
  inv1 g18627(.a(new_n18808), .O(new_n18821));
  inv1 g18628(.a(new_n18819), .O(new_n18822));
  nor2 g18629(.a(new_n18822), .b(new_n18821), .O(new_n18823));
  nor2 g18630(.a(new_n18823), .b(new_n18820), .O(new_n18824));
  nor2 g18631(.a(new_n18824), .b(new_n18795), .O(new_n18825));
  inv1 g18632(.a(new_n18824), .O(new_n18826));
  nor2 g18633(.a(new_n18826), .b(new_n18794), .O(new_n18827));
  nor2 g18634(.a(new_n18827), .b(new_n18825), .O(new_n18828));
  nor2 g18635(.a(new_n18828), .b(new_n18781), .O(new_n18829));
  inv1 g18636(.a(new_n18781), .O(new_n18830));
  inv1 g18637(.a(new_n18828), .O(new_n18831));
  nor2 g18638(.a(new_n18831), .b(new_n18830), .O(new_n18832));
  nor2 g18639(.a(new_n18832), .b(new_n18829), .O(new_n18833));
  inv1 g18640(.a(new_n18833), .O(new_n18834));
  nor2 g18641(.a(new_n9873), .b(new_n2506), .O(new_n18835));
  nor2 g18642(.a(new_n7537), .b(new_n3870), .O(new_n18836));
  nor2 g18643(.a(new_n18836), .b(new_n18835), .O(new_n18837));
  inv1 g18644(.a(new_n18835), .O(new_n18838));
  inv1 g18645(.a(new_n18836), .O(new_n18839));
  nor2 g18646(.a(new_n18839), .b(new_n18838), .O(new_n18840));
  nor2 g18647(.a(new_n18840), .b(new_n18837), .O(new_n18841));
  nor2 g18648(.a(new_n18841), .b(new_n18670), .O(new_n18842));
  inv1 g18649(.a(new_n18841), .O(new_n18843));
  nor2 g18650(.a(new_n18843), .b(new_n18669), .O(new_n18844));
  nor2 g18651(.a(new_n18844), .b(new_n18842), .O(new_n18845));
  nor2 g18652(.a(new_n8170), .b(new_n3533), .O(new_n18846));
  nor2 g18653(.a(new_n18846), .b(new_n18170), .O(new_n18847));
  inv1 g18654(.a(new_n18846), .O(new_n18848));
  nor2 g18655(.a(new_n18848), .b(new_n18171), .O(new_n18849));
  nor2 g18656(.a(new_n18849), .b(new_n18847), .O(new_n18850));
  nor2 g18657(.a(new_n18850), .b(new_n18611), .O(new_n18851));
  inv1 g18658(.a(new_n18850), .O(new_n18852));
  nor2 g18659(.a(new_n18852), .b(new_n18610), .O(new_n18853));
  nor2 g18660(.a(new_n18853), .b(new_n18851), .O(new_n18854));
  nor2 g18661(.a(new_n18506), .b(new_n18501), .O(new_n18855));
  nor2 g18662(.a(new_n18855), .b(new_n18854), .O(new_n18856));
  inv1 g18663(.a(new_n18854), .O(new_n18857));
  inv1 g18664(.a(new_n18855), .O(new_n18858));
  nor2 g18665(.a(new_n18858), .b(new_n18857), .O(new_n18859));
  nor2 g18666(.a(new_n18859), .b(new_n18856), .O(new_n18860));
  inv1 g18667(.a(new_n18860), .O(new_n18861));
  nor2 g18668(.a(new_n18861), .b(new_n18845), .O(new_n18862));
  inv1 g18669(.a(new_n18845), .O(new_n18863));
  nor2 g18670(.a(new_n18860), .b(new_n18863), .O(new_n18864));
  nor2 g18671(.a(new_n18864), .b(new_n18862), .O(new_n18865));
  inv1 g18672(.a(new_n18865), .O(new_n18866));
  nor2 g18673(.a(new_n18866), .b(new_n18834), .O(new_n18867));
  nor2 g18674(.a(new_n18865), .b(new_n18833), .O(new_n18868));
  nor2 g18675(.a(new_n18868), .b(new_n18867), .O(new_n18869));
  inv1 g18676(.a(new_n18869), .O(new_n18870));
  nor2 g18677(.a(new_n18870), .b(new_n18753), .O(new_n18871));
  inv1 g18678(.a(new_n18753), .O(new_n18872));
  nor2 g18679(.a(new_n18869), .b(new_n18872), .O(new_n18873));
  nor2 g18680(.a(new_n18873), .b(new_n18871), .O(new_n18874));
  inv1 g18681(.a(new_n18874), .O(new_n18875));
  nor2 g18682(.a(new_n18583), .b(new_n18579), .O(new_n18876));
  inv1 g18683(.a(new_n18876), .O(new_n18877));
  nor2 g18684(.a(new_n18547), .b(new_n18541), .O(new_n18878));
  inv1 g18685(.a(new_n18878), .O(new_n18879));
  nor2 g18686(.a(new_n18879), .b(new_n18877), .O(new_n18880));
  nor2 g18687(.a(new_n18878), .b(new_n18876), .O(new_n18881));
  nor2 g18688(.a(new_n18881), .b(new_n18880), .O(new_n18882));
  inv1 g18689(.a(new_n18882), .O(new_n18883));
  nor2 g18690(.a(new_n18517), .b(new_n18511), .O(new_n18884));
  nor2 g18691(.a(new_n18628), .b(new_n18621), .O(new_n18885));
  nor2 g18692(.a(new_n18604), .b(new_n18597), .O(new_n18886));
  nor2 g18693(.a(new_n18886), .b(new_n18885), .O(new_n18887));
  inv1 g18694(.a(new_n18885), .O(new_n18888));
  inv1 g18695(.a(new_n18886), .O(new_n18889));
  nor2 g18696(.a(new_n18889), .b(new_n18888), .O(new_n18890));
  nor2 g18697(.a(new_n18890), .b(new_n18887), .O(new_n18891));
  nor2 g18698(.a(new_n18648), .b(new_n18641), .O(new_n18892));
  nor2 g18699(.a(new_n18892), .b(new_n18891), .O(new_n18893));
  inv1 g18700(.a(new_n18891), .O(new_n18894));
  inv1 g18701(.a(new_n18892), .O(new_n18895));
  nor2 g18702(.a(new_n18895), .b(new_n18894), .O(new_n18896));
  nor2 g18703(.a(new_n18896), .b(new_n18893), .O(new_n18897));
  nor2 g18704(.a(new_n18675), .b(new_n18667), .O(new_n18898));
  nor2 g18705(.a(new_n18615), .b(new_n18608), .O(new_n18899));
  nor2 g18706(.a(new_n18899), .b(new_n18898), .O(new_n18900));
  inv1 g18707(.a(new_n18898), .O(new_n18901));
  inv1 g18708(.a(new_n18899), .O(new_n18902));
  nor2 g18709(.a(new_n18902), .b(new_n18901), .O(new_n18903));
  nor2 g18710(.a(new_n18903), .b(new_n18900), .O(new_n18904));
  nor2 g18711(.a(new_n18660), .b(new_n18654), .O(new_n18905));
  nor2 g18712(.a(new_n18905), .b(new_n18904), .O(new_n18906));
  inv1 g18713(.a(new_n18904), .O(new_n18907));
  inv1 g18714(.a(new_n18905), .O(new_n18908));
  nor2 g18715(.a(new_n18908), .b(new_n18907), .O(new_n18909));
  nor2 g18716(.a(new_n18909), .b(new_n18906), .O(new_n18910));
  nor2 g18717(.a(new_n18910), .b(new_n18897), .O(new_n18911));
  inv1 g18718(.a(new_n18897), .O(new_n18912));
  inv1 g18719(.a(new_n18910), .O(new_n18913));
  nor2 g18720(.a(new_n18913), .b(new_n18912), .O(new_n18914));
  nor2 g18721(.a(new_n18914), .b(new_n18911), .O(new_n18915));
  inv1 g18722(.a(new_n18915), .O(new_n18916));
  nor2 g18723(.a(new_n18916), .b(new_n18884), .O(new_n18917));
  inv1 g18724(.a(new_n18884), .O(new_n18918));
  nor2 g18725(.a(new_n18915), .b(new_n18918), .O(new_n18919));
  nor2 g18726(.a(new_n18919), .b(new_n18917), .O(new_n18920));
  inv1 g18727(.a(new_n18920), .O(new_n18921));
  nor2 g18728(.a(new_n18921), .b(new_n18883), .O(new_n18922));
  nor2 g18729(.a(new_n18920), .b(new_n18882), .O(new_n18923));
  nor2 g18730(.a(new_n18923), .b(new_n18922), .O(new_n18924));
  inv1 g18731(.a(new_n18924), .O(new_n18925));
  nor2 g18732(.a(new_n18925), .b(new_n18875), .O(new_n18926));
  nor2 g18733(.a(new_n18924), .b(new_n18874), .O(new_n18927));
  nor2 g18734(.a(new_n18927), .b(new_n18926), .O(new_n18928));
  nor2 g18735(.a(new_n18928), .b(new_n18752), .O(new_n18929));
  inv1 g18736(.a(new_n18752), .O(new_n18930));
  inv1 g18737(.a(new_n18928), .O(new_n18931));
  nor2 g18738(.a(new_n18931), .b(new_n18930), .O(new_n18932));
  nor2 g18739(.a(new_n18932), .b(new_n18929), .O(new_n18933));
  nor2 g18740(.a(new_n18933), .b(new_n18721), .O(new_n18934));
  inv1 g18741(.a(new_n18933), .O(new_n18935));
  nor2 g18742(.a(new_n18935), .b(new_n18720), .O(new_n18936));
  nor2 g18743(.a(new_n18936), .b(new_n18934), .O(new_n18937));
  inv1 g18744(.a(new_n18937), .O(new_n18938));
  nor2 g18745(.a(new_n18717), .b(new_n18709), .O(new_n18939));
  nor2 g18746(.a(new_n18939), .b(new_n18938), .O(new_n18940));
  inv1 g18747(.a(new_n18939), .O(new_n18941));
  nor2 g18748(.a(new_n18941), .b(new_n18937), .O(new_n18942));
  nor2 g18749(.a(new_n18942), .b(new_n18940), .O(new_n18943));
  inv1 g18750(.a(new_n18943), .O(\asquared[88] ));
  nor2 g18751(.a(new_n18932), .b(new_n18751), .O(new_n18945));
  inv1 g18752(.a(new_n18945), .O(new_n18946));
  nor2 g18753(.a(new_n18926), .b(new_n18871), .O(new_n18947));
  nor2 g18754(.a(new_n18922), .b(new_n18881), .O(new_n18948));
  nor2 g18755(.a(new_n18909), .b(new_n18903), .O(new_n18949));
  inv1 g18756(.a(new_n18949), .O(new_n18950));
  nor2 g18757(.a(new_n18862), .b(new_n18856), .O(new_n18951));
  inv1 g18758(.a(new_n18951), .O(new_n18952));
  nor2 g18759(.a(new_n18952), .b(new_n18950), .O(new_n18953));
  nor2 g18760(.a(new_n18951), .b(new_n18949), .O(new_n18954));
  nor2 g18761(.a(new_n18954), .b(new_n18953), .O(new_n18955));
  nor2 g18762(.a(new_n18827), .b(new_n18820), .O(new_n18956));
  inv1 g18763(.a(new_n18956), .O(new_n18957));
  nor2 g18764(.a(new_n18957), .b(new_n18955), .O(new_n18958));
  inv1 g18765(.a(new_n18955), .O(new_n18959));
  nor2 g18766(.a(new_n18956), .b(new_n18959), .O(new_n18960));
  nor2 g18767(.a(new_n18960), .b(new_n18958), .O(new_n18961));
  inv1 g18768(.a(new_n18961), .O(new_n18962));
  nor2 g18769(.a(new_n18867), .b(new_n18832), .O(new_n18963));
  nor2 g18770(.a(new_n18963), .b(new_n18962), .O(new_n18964));
  inv1 g18771(.a(new_n18963), .O(new_n18965));
  nor2 g18772(.a(new_n18965), .b(new_n18961), .O(new_n18966));
  nor2 g18773(.a(new_n18966), .b(new_n18964), .O(new_n18967));
  inv1 g18774(.a(new_n18967), .O(new_n18968));
  nor2 g18775(.a(new_n18968), .b(new_n18948), .O(new_n18969));
  inv1 g18776(.a(new_n18948), .O(new_n18970));
  nor2 g18777(.a(new_n18967), .b(new_n18970), .O(new_n18971));
  nor2 g18778(.a(new_n18971), .b(new_n18969), .O(new_n18972));
  inv1 g18779(.a(new_n18972), .O(new_n18973));
  nor2 g18780(.a(new_n18973), .b(new_n18947), .O(new_n18974));
  inv1 g18781(.a(new_n18947), .O(new_n18975));
  nor2 g18782(.a(new_n18972), .b(new_n18975), .O(new_n18976));
  nor2 g18783(.a(new_n18976), .b(new_n18974), .O(new_n18977));
  nor2 g18784(.a(new_n18917), .b(new_n18914), .O(new_n18978));
  inv1 g18785(.a(new_n18978), .O(new_n18979));
  nor2 g18786(.a(new_n18734), .b(new_n18728), .O(new_n18980));
  inv1 g18787(.a(new_n18980), .O(new_n18981));
  nor2 g18788(.a(new_n18981), .b(new_n18979), .O(new_n18982));
  nor2 g18789(.a(new_n18980), .b(new_n18978), .O(new_n18983));
  nor2 g18790(.a(new_n18983), .b(new_n18982), .O(new_n18984));
  inv1 g18791(.a(new_n18984), .O(new_n18985));
  nor2 g18792(.a(new_n18853), .b(new_n18847), .O(new_n18986));
  nor2 g18793(.a(new_n18805), .b(new_n18799), .O(new_n18987));
  nor2 g18794(.a(new_n18987), .b(new_n18986), .O(new_n18988));
  inv1 g18795(.a(new_n18986), .O(new_n18989));
  inv1 g18796(.a(new_n18987), .O(new_n18990));
  nor2 g18797(.a(new_n18990), .b(new_n18989), .O(new_n18991));
  nor2 g18798(.a(new_n18991), .b(new_n18988), .O(new_n18992));
  nor2 g18799(.a(new_n18818), .b(new_n18811), .O(new_n18993));
  nor2 g18800(.a(new_n18993), .b(new_n18992), .O(new_n18994));
  inv1 g18801(.a(new_n18992), .O(new_n18995));
  inv1 g18802(.a(new_n18993), .O(new_n18996));
  nor2 g18803(.a(new_n18996), .b(new_n18995), .O(new_n18997));
  nor2 g18804(.a(new_n18997), .b(new_n18994), .O(new_n18998));
  inv1 g18805(.a(new_n18998), .O(new_n18999));
  nor2 g18806(.a(new_n18780), .b(new_n18773), .O(new_n19000));
  inv1 g18807(.a(new_n19000), .O(new_n19001));
  nor2 g18808(.a(new_n18844), .b(new_n18837), .O(new_n19002));
  nor2 g18809(.a(new_n18766), .b(new_n18758), .O(new_n19003));
  nor2 g18810(.a(new_n19003), .b(new_n19002), .O(new_n19004));
  inv1 g18811(.a(new_n19002), .O(new_n19005));
  inv1 g18812(.a(new_n19003), .O(new_n19006));
  nor2 g18813(.a(new_n19006), .b(new_n19005), .O(new_n19007));
  nor2 g18814(.a(new_n19007), .b(new_n19004), .O(new_n19008));
  inv1 g18815(.a(new_n19008), .O(new_n19009));
  nor2 g18816(.a(new_n5971), .b(new_n5393), .O(new_n19010));
  inv1 g18817(.a(new_n19010), .O(new_n19011));
  nor2 g18818(.a(new_n8946), .b(new_n3231), .O(new_n19012));
  nor2 g18819(.a(new_n8476), .b(new_n3533), .O(new_n19013));
  nor2 g18820(.a(new_n19013), .b(new_n19012), .O(new_n19014));
  inv1 g18821(.a(new_n18757), .O(new_n19015));
  nor2 g18822(.a(new_n8946), .b(new_n3533), .O(new_n19016));
  inv1 g18823(.a(new_n19016), .O(new_n19017));
  nor2 g18824(.a(new_n19017), .b(new_n19015), .O(new_n19018));
  nor2 g18825(.a(new_n19018), .b(new_n19014), .O(new_n19019));
  nor2 g18826(.a(new_n19019), .b(new_n19011), .O(new_n19020));
  inv1 g18827(.a(new_n19019), .O(new_n19021));
  nor2 g18828(.a(new_n19021), .b(new_n19010), .O(new_n19022));
  nor2 g18829(.a(new_n19022), .b(new_n19020), .O(new_n19023));
  nor2 g18830(.a(new_n19023), .b(new_n19009), .O(new_n19024));
  inv1 g18831(.a(new_n19023), .O(new_n19025));
  nor2 g18832(.a(new_n19025), .b(new_n19008), .O(new_n19026));
  nor2 g18833(.a(new_n19026), .b(new_n19024), .O(new_n19027));
  nor2 g18834(.a(new_n19027), .b(new_n19001), .O(new_n19028));
  inv1 g18835(.a(new_n19027), .O(new_n19029));
  nor2 g18836(.a(new_n19029), .b(new_n19000), .O(new_n19030));
  nor2 g18837(.a(new_n19030), .b(new_n19028), .O(new_n19031));
  inv1 g18838(.a(new_n19031), .O(new_n19032));
  nor2 g18839(.a(new_n19032), .b(new_n18999), .O(new_n19033));
  nor2 g18840(.a(new_n19031), .b(new_n18998), .O(new_n19034));
  nor2 g18841(.a(new_n19034), .b(new_n19033), .O(new_n19035));
  inv1 g18842(.a(new_n19035), .O(new_n19036));
  nor2 g18843(.a(new_n19036), .b(new_n18985), .O(new_n19037));
  nor2 g18844(.a(new_n19035), .b(new_n18984), .O(new_n19038));
  nor2 g18845(.a(new_n19038), .b(new_n19037), .O(new_n19039));
  inv1 g18846(.a(new_n19039), .O(new_n19040));
  nor2 g18847(.a(new_n18745), .b(new_n18737), .O(new_n19041));
  nor2 g18848(.a(new_n18896), .b(new_n18890), .O(new_n19042));
  inv1 g18849(.a(new_n19042), .O(new_n19043));
  nor2 g18850(.a(new_n10320), .b(new_n2506), .O(new_n19044));
  nor2 g18851(.a(new_n7294), .b(new_n4366), .O(new_n19045));
  nor2 g18852(.a(new_n19045), .b(new_n18812), .O(new_n19046));
  inv1 g18853(.a(new_n18809), .O(new_n19047));
  nor2 g18854(.a(new_n7294), .b(new_n4425), .O(new_n19048));
  inv1 g18855(.a(new_n19048), .O(new_n19049));
  nor2 g18856(.a(new_n19049), .b(new_n19047), .O(new_n19050));
  nor2 g18857(.a(new_n19050), .b(new_n19046), .O(new_n19051));
  inv1 g18858(.a(new_n19051), .O(new_n19052));
  nor2 g18859(.a(new_n19052), .b(new_n19044), .O(new_n19053));
  inv1 g18860(.a(new_n19044), .O(new_n19054));
  nor2 g18861(.a(new_n19051), .b(new_n19054), .O(new_n19055));
  nor2 g18862(.a(new_n19055), .b(new_n19053), .O(new_n19056));
  nor2 g18863(.a(new_n6893), .b(new_n4682), .O(new_n19057));
  inv1 g18864(.a(new_n19057), .O(new_n19058));
  nor2 g18865(.a(new_n9873), .b(new_n2660), .O(new_n19059));
  nor2 g18866(.a(new_n9156), .b(new_n3057), .O(new_n19060));
  nor2 g18867(.a(new_n19060), .b(new_n19059), .O(new_n19061));
  nor2 g18868(.a(new_n9873), .b(new_n3057), .O(new_n19062));
  inv1 g18869(.a(new_n19062), .O(new_n19063));
  nor2 g18870(.a(new_n19063), .b(new_n18594), .O(new_n19064));
  nor2 g18871(.a(new_n19064), .b(new_n19061), .O(new_n19065));
  nor2 g18872(.a(new_n19065), .b(new_n19058), .O(new_n19066));
  inv1 g18873(.a(new_n19065), .O(new_n19067));
  nor2 g18874(.a(new_n19067), .b(new_n19057), .O(new_n19068));
  nor2 g18875(.a(new_n19068), .b(new_n19066), .O(new_n19069));
  nor2 g18876(.a(new_n19069), .b(new_n19056), .O(new_n19070));
  inv1 g18877(.a(new_n19056), .O(new_n19071));
  inv1 g18878(.a(new_n19069), .O(new_n19072));
  nor2 g18879(.a(new_n19072), .b(new_n19071), .O(new_n19073));
  nor2 g18880(.a(new_n19073), .b(new_n19070), .O(new_n19074));
  nor2 g18881(.a(new_n19074), .b(new_n19043), .O(new_n19075));
  inv1 g18882(.a(new_n19074), .O(new_n19076));
  nor2 g18883(.a(new_n19076), .b(new_n19042), .O(new_n19077));
  nor2 g18884(.a(new_n19077), .b(new_n19075), .O(new_n19078));
  inv1 g18885(.a(new_n19078), .O(new_n19079));
  nor2 g18886(.a(new_n11596), .b(new_n1903), .O(new_n19080));
  inv1 g18887(.a(new_n19080), .O(new_n19081));
  nor2 g18888(.a(new_n18771), .b(new_n5796), .O(new_n19082));
  inv1 g18889(.a(new_n19082), .O(new_n19083));
  nor2 g18890(.a(new_n19083), .b(new_n19081), .O(new_n19084));
  nor2 g18891(.a(new_n19082), .b(new_n19080), .O(new_n19085));
  nor2 g18892(.a(new_n19085), .b(new_n19084), .O(new_n19086));
  nor2 g18893(.a(new_n18793), .b(new_n18786), .O(new_n19087));
  nor2 g18894(.a(new_n19087), .b(new_n19086), .O(new_n19088));
  inv1 g18895(.a(new_n19086), .O(new_n19089));
  inv1 g18896(.a(new_n19087), .O(new_n19090));
  nor2 g18897(.a(new_n19090), .b(new_n19089), .O(new_n19091));
  nor2 g18898(.a(new_n19091), .b(new_n19088), .O(new_n19092));
  inv1 g18899(.a(new_n19092), .O(new_n19093));
  nor2 g18900(.a(new_n19093), .b(new_n19079), .O(new_n19094));
  nor2 g18901(.a(new_n19092), .b(new_n19078), .O(new_n19095));
  nor2 g18902(.a(new_n19095), .b(new_n19094), .O(new_n19096));
  inv1 g18903(.a(new_n19096), .O(new_n19097));
  nor2 g18904(.a(new_n8170), .b(new_n3722), .O(new_n19098));
  inv1 g18905(.a(new_n19098), .O(new_n19099));
  nor2 g18906(.a(new_n7537), .b(new_n4093), .O(new_n19100));
  nor2 g18907(.a(new_n8026), .b(new_n3870), .O(new_n19101));
  nor2 g18908(.a(new_n19101), .b(new_n19100), .O(new_n19102));
  nor2 g18909(.a(new_n8026), .b(new_n4093), .O(new_n19103));
  inv1 g18910(.a(new_n19103), .O(new_n19104));
  nor2 g18911(.a(new_n19104), .b(new_n18839), .O(new_n19105));
  nor2 g18912(.a(new_n19105), .b(new_n19102), .O(new_n19106));
  nor2 g18913(.a(new_n19106), .b(new_n19099), .O(new_n19107));
  inv1 g18914(.a(new_n19106), .O(new_n19108));
  nor2 g18915(.a(new_n19108), .b(new_n19098), .O(new_n19109));
  nor2 g18916(.a(new_n19109), .b(new_n19107), .O(new_n19110));
  inv1 g18917(.a(new_n19110), .O(new_n19111));
  nor2 g18918(.a(new_n11186), .b(new_n2121), .O(new_n19112));
  nor2 g18919(.a(new_n10468), .b(new_n2433), .O(new_n19113));
  nor2 g18920(.a(new_n19113), .b(new_n18800), .O(new_n19114));
  inv1 g18921(.a(new_n18798), .O(new_n19115));
  nor2 g18922(.a(new_n10895), .b(new_n2433), .O(new_n19116));
  inv1 g18923(.a(new_n19116), .O(new_n19117));
  nor2 g18924(.a(new_n19117), .b(new_n19115), .O(new_n19118));
  nor2 g18925(.a(new_n19118), .b(new_n19114), .O(new_n19119));
  inv1 g18926(.a(new_n19119), .O(new_n19120));
  nor2 g18927(.a(new_n19120), .b(new_n19112), .O(new_n19121));
  inv1 g18928(.a(new_n19112), .O(new_n19122));
  nor2 g18929(.a(new_n19119), .b(new_n19122), .O(new_n19123));
  nor2 g18930(.a(new_n19123), .b(new_n19121), .O(new_n19124));
  nor2 g18931(.a(new_n6570), .b(new_n4954), .O(new_n19125));
  nor2 g18932(.a(new_n19125), .b(new_n18787), .O(new_n19126));
  inv1 g18933(.a(new_n18785), .O(new_n19127));
  nor2 g18934(.a(new_n6570), .b(new_n5178), .O(new_n19128));
  inv1 g18935(.a(new_n19128), .O(new_n19129));
  nor2 g18936(.a(new_n19129), .b(new_n19127), .O(new_n19130));
  nor2 g18937(.a(new_n19130), .b(new_n19126), .O(new_n19131));
  nor2 g18938(.a(new_n19131), .b(new_n18643), .O(new_n19132));
  inv1 g18939(.a(new_n19131), .O(new_n19133));
  nor2 g18940(.a(new_n19133), .b(new_n18642), .O(new_n19134));
  nor2 g18941(.a(new_n19134), .b(new_n19132), .O(new_n19135));
  nor2 g18942(.a(new_n19135), .b(new_n19124), .O(new_n19136));
  inv1 g18943(.a(new_n19124), .O(new_n19137));
  inv1 g18944(.a(new_n19135), .O(new_n19138));
  nor2 g18945(.a(new_n19138), .b(new_n19137), .O(new_n19139));
  nor2 g18946(.a(new_n19139), .b(new_n19136), .O(new_n19140));
  nor2 g18947(.a(new_n19140), .b(new_n19111), .O(new_n19141));
  inv1 g18948(.a(new_n19140), .O(new_n19142));
  nor2 g18949(.a(new_n19142), .b(new_n19110), .O(new_n19143));
  nor2 g18950(.a(new_n19143), .b(new_n19141), .O(new_n19144));
  inv1 g18951(.a(new_n19144), .O(new_n19145));
  nor2 g18952(.a(new_n19145), .b(new_n19097), .O(new_n19146));
  nor2 g18953(.a(new_n19144), .b(new_n19096), .O(new_n19147));
  nor2 g18954(.a(new_n19147), .b(new_n19146), .O(new_n19148));
  inv1 g18955(.a(new_n19148), .O(new_n19149));
  nor2 g18956(.a(new_n19149), .b(new_n19041), .O(new_n19150));
  inv1 g18957(.a(new_n19041), .O(new_n19151));
  nor2 g18958(.a(new_n19148), .b(new_n19151), .O(new_n19152));
  nor2 g18959(.a(new_n19152), .b(new_n19150), .O(new_n19153));
  inv1 g18960(.a(new_n19153), .O(new_n19154));
  nor2 g18961(.a(new_n19154), .b(new_n19040), .O(new_n19155));
  nor2 g18962(.a(new_n19153), .b(new_n19039), .O(new_n19156));
  nor2 g18963(.a(new_n19156), .b(new_n19155), .O(new_n19157));
  inv1 g18964(.a(new_n19157), .O(new_n19158));
  nor2 g18965(.a(new_n19158), .b(new_n18977), .O(new_n19159));
  inv1 g18966(.a(new_n18977), .O(new_n19160));
  nor2 g18967(.a(new_n19157), .b(new_n19160), .O(new_n19161));
  nor2 g18968(.a(new_n19161), .b(new_n19159), .O(new_n19162));
  inv1 g18969(.a(new_n19162), .O(new_n19163));
  nor2 g18970(.a(new_n19163), .b(new_n18946), .O(new_n19164));
  nor2 g18971(.a(new_n19162), .b(new_n18945), .O(new_n19165));
  nor2 g18972(.a(new_n19165), .b(new_n19164), .O(new_n19166));
  inv1 g18973(.a(new_n19166), .O(new_n19167));
  nor2 g18974(.a(new_n18940), .b(new_n18934), .O(new_n19168));
  inv1 g18975(.a(new_n19168), .O(new_n19169));
  nor2 g18976(.a(new_n19169), .b(new_n19167), .O(new_n19170));
  nor2 g18977(.a(new_n19168), .b(new_n19166), .O(new_n19171));
  nor2 g18978(.a(new_n19171), .b(new_n19170), .O(\asquared[89] ));
  nor2 g18979(.a(new_n18997), .b(new_n18991), .O(new_n19173));
  inv1 g18980(.a(new_n19173), .O(new_n19174));
  nor2 g18981(.a(new_n19091), .b(new_n19084), .O(new_n19175));
  inv1 g18982(.a(new_n19175), .O(new_n19176));
  nor2 g18983(.a(new_n19176), .b(new_n19174), .O(new_n19177));
  nor2 g18984(.a(new_n19175), .b(new_n19173), .O(new_n19178));
  nor2 g18985(.a(new_n19178), .b(new_n19177), .O(new_n19179));
  nor2 g18986(.a(new_n19024), .b(new_n19007), .O(new_n19180));
  inv1 g18987(.a(new_n19180), .O(new_n19181));
  nor2 g18988(.a(new_n19181), .b(new_n19179), .O(new_n19182));
  inv1 g18989(.a(new_n19179), .O(new_n19183));
  nor2 g18990(.a(new_n19180), .b(new_n19183), .O(new_n19184));
  nor2 g18991(.a(new_n19184), .b(new_n19182), .O(new_n19185));
  nor2 g18992(.a(new_n18960), .b(new_n18954), .O(new_n19186));
  inv1 g18993(.a(new_n19186), .O(new_n19187));
  nor2 g18994(.a(new_n19187), .b(new_n19185), .O(new_n19188));
  inv1 g18995(.a(new_n19185), .O(new_n19189));
  nor2 g18996(.a(new_n19186), .b(new_n19189), .O(new_n19190));
  nor2 g18997(.a(new_n19190), .b(new_n19188), .O(new_n19191));
  inv1 g18998(.a(new_n19191), .O(new_n19192));
  nor2 g18999(.a(new_n19033), .b(new_n19030), .O(new_n19193));
  nor2 g19000(.a(new_n19193), .b(new_n19192), .O(new_n19194));
  inv1 g19001(.a(new_n19193), .O(new_n19195));
  nor2 g19002(.a(new_n19195), .b(new_n19191), .O(new_n19196));
  nor2 g19003(.a(new_n19196), .b(new_n19194), .O(new_n19197));
  inv1 g19004(.a(new_n19197), .O(new_n19198));
  nor2 g19005(.a(new_n18969), .b(new_n18964), .O(new_n19199));
  nor2 g19006(.a(new_n19109), .b(new_n19102), .O(new_n19200));
  nor2 g19007(.a(new_n19121), .b(new_n19114), .O(new_n19201));
  nor2 g19008(.a(new_n19201), .b(new_n19200), .O(new_n19202));
  inv1 g19009(.a(new_n19200), .O(new_n19203));
  inv1 g19010(.a(new_n19201), .O(new_n19204));
  nor2 g19011(.a(new_n19204), .b(new_n19203), .O(new_n19205));
  nor2 g19012(.a(new_n19205), .b(new_n19202), .O(new_n19206));
  nor2 g19013(.a(new_n19068), .b(new_n19061), .O(new_n19207));
  nor2 g19014(.a(new_n19207), .b(new_n19206), .O(new_n19208));
  inv1 g19015(.a(new_n19206), .O(new_n19209));
  inv1 g19016(.a(new_n19207), .O(new_n19210));
  nor2 g19017(.a(new_n19210), .b(new_n19209), .O(new_n19211));
  nor2 g19018(.a(new_n19211), .b(new_n19208), .O(new_n19212));
  inv1 g19019(.a(new_n19212), .O(new_n19213));
  nor2 g19020(.a(new_n10468), .b(new_n2506), .O(new_n19214));
  nor2 g19021(.a(new_n19214), .b(new_n19116), .O(new_n19215));
  inv1 g19022(.a(new_n19113), .O(new_n19216));
  nor2 g19023(.a(new_n10895), .b(new_n2506), .O(new_n19217));
  inv1 g19024(.a(new_n19217), .O(new_n19218));
  nor2 g19025(.a(new_n19218), .b(new_n19216), .O(new_n19219));
  nor2 g19026(.a(new_n19219), .b(new_n19215), .O(new_n19220));
  inv1 g19027(.a(new_n19220), .O(new_n19221));
  nor2 g19028(.a(new_n19022), .b(new_n19014), .O(new_n19222));
  inv1 g19029(.a(new_n19222), .O(new_n19223));
  nor2 g19030(.a(new_n19223), .b(new_n19221), .O(new_n19224));
  nor2 g19031(.a(new_n19222), .b(new_n19220), .O(new_n19225));
  nor2 g19032(.a(new_n19225), .b(new_n19224), .O(new_n19226));
  inv1 g19033(.a(new_n19226), .O(new_n19227));
  nor2 g19034(.a(new_n6274), .b(new_n5393), .O(new_n19228));
  nor2 g19035(.a(new_n19228), .b(new_n19128), .O(new_n19229));
  nor2 g19036(.a(new_n6570), .b(new_n5393), .O(new_n19230));
  inv1 g19037(.a(new_n19230), .O(new_n19231));
  nor2 g19038(.a(new_n19231), .b(new_n18788), .O(new_n19232));
  nor2 g19039(.a(new_n19232), .b(new_n19229), .O(new_n19233));
  nor2 g19040(.a(new_n19233), .b(new_n19017), .O(new_n19234));
  inv1 g19041(.a(new_n19233), .O(new_n19235));
  nor2 g19042(.a(new_n19235), .b(new_n19016), .O(new_n19236));
  nor2 g19043(.a(new_n19236), .b(new_n19234), .O(new_n19237));
  nor2 g19044(.a(new_n11186), .b(new_n2184), .O(new_n19238));
  inv1 g19045(.a(new_n19238), .O(new_n19239));
  nor2 g19046(.a(new_n5971), .b(\a[44] ), .O(new_n19240));
  nor2 g19047(.a(new_n19240), .b(new_n19239), .O(new_n19241));
  inv1 g19048(.a(new_n19240), .O(new_n19242));
  nor2 g19049(.a(new_n19242), .b(new_n19238), .O(new_n19243));
  nor2 g19050(.a(new_n19243), .b(new_n19241), .O(new_n19244));
  nor2 g19051(.a(new_n19244), .b(new_n19237), .O(new_n19245));
  inv1 g19052(.a(new_n19237), .O(new_n19246));
  inv1 g19053(.a(new_n19244), .O(new_n19247));
  nor2 g19054(.a(new_n19247), .b(new_n19246), .O(new_n19248));
  nor2 g19055(.a(new_n19248), .b(new_n19245), .O(new_n19249));
  inv1 g19056(.a(new_n19249), .O(new_n19250));
  nor2 g19057(.a(new_n19250), .b(new_n19227), .O(new_n19251));
  nor2 g19058(.a(new_n19249), .b(new_n19226), .O(new_n19252));
  nor2 g19059(.a(new_n19252), .b(new_n19251), .O(new_n19253));
  inv1 g19060(.a(new_n19253), .O(new_n19254));
  nor2 g19061(.a(new_n19254), .b(new_n19213), .O(new_n19255));
  nor2 g19062(.a(new_n19253), .b(new_n19212), .O(new_n19256));
  nor2 g19063(.a(new_n19256), .b(new_n19255), .O(new_n19257));
  inv1 g19064(.a(new_n19257), .O(new_n19258));
  nor2 g19065(.a(new_n10320), .b(new_n2660), .O(new_n19259));
  inv1 g19066(.a(new_n19259), .O(new_n19260));
  nor2 g19067(.a(new_n9873), .b(new_n2826), .O(new_n19261));
  nor2 g19068(.a(new_n19261), .b(new_n17810), .O(new_n19262));
  nor2 g19069(.a(new_n19063), .b(new_n18643), .O(new_n19263));
  nor2 g19070(.a(new_n19263), .b(new_n19262), .O(new_n19264));
  nor2 g19071(.a(new_n19264), .b(new_n19260), .O(new_n19265));
  inv1 g19072(.a(new_n19264), .O(new_n19266));
  nor2 g19073(.a(new_n19266), .b(new_n19259), .O(new_n19267));
  nor2 g19074(.a(new_n19267), .b(new_n19265), .O(new_n19268));
  inv1 g19075(.a(new_n19268), .O(new_n19269));
  nor2 g19076(.a(new_n6893), .b(new_n4954), .O(new_n19270));
  nor2 g19077(.a(new_n8476), .b(new_n3722), .O(new_n19271));
  nor2 g19078(.a(new_n19271), .b(new_n18760), .O(new_n19272));
  nor2 g19079(.a(new_n9156), .b(new_n3722), .O(new_n19273));
  inv1 g19080(.a(new_n19273), .O(new_n19274));
  nor2 g19081(.a(new_n19274), .b(new_n19015), .O(new_n19275));
  nor2 g19082(.a(new_n19275), .b(new_n19272), .O(new_n19276));
  inv1 g19083(.a(new_n19276), .O(new_n19277));
  nor2 g19084(.a(new_n19277), .b(new_n19270), .O(new_n19278));
  inv1 g19085(.a(new_n19270), .O(new_n19279));
  nor2 g19086(.a(new_n19276), .b(new_n19279), .O(new_n19280));
  nor2 g19087(.a(new_n19280), .b(new_n19278), .O(new_n19281));
  nor2 g19088(.a(new_n8170), .b(new_n3870), .O(new_n19282));
  inv1 g19089(.a(new_n19282), .O(new_n19283));
  nor2 g19090(.a(new_n7537), .b(new_n4366), .O(new_n19284));
  nor2 g19091(.a(new_n19284), .b(new_n19103), .O(new_n19285));
  inv1 g19092(.a(new_n19100), .O(new_n19286));
  nor2 g19093(.a(new_n8026), .b(new_n4366), .O(new_n19287));
  inv1 g19094(.a(new_n19287), .O(new_n19288));
  nor2 g19095(.a(new_n19288), .b(new_n19286), .O(new_n19289));
  nor2 g19096(.a(new_n19289), .b(new_n19285), .O(new_n19290));
  nor2 g19097(.a(new_n19290), .b(new_n19283), .O(new_n19291));
  inv1 g19098(.a(new_n19290), .O(new_n19292));
  nor2 g19099(.a(new_n19292), .b(new_n19282), .O(new_n19293));
  nor2 g19100(.a(new_n19293), .b(new_n19291), .O(new_n19294));
  nor2 g19101(.a(new_n19294), .b(new_n19281), .O(new_n19295));
  inv1 g19102(.a(new_n19281), .O(new_n19296));
  inv1 g19103(.a(new_n19294), .O(new_n19297));
  nor2 g19104(.a(new_n19297), .b(new_n19296), .O(new_n19298));
  nor2 g19105(.a(new_n19298), .b(new_n19295), .O(new_n19299));
  nor2 g19106(.a(new_n19299), .b(new_n19269), .O(new_n19300));
  inv1 g19107(.a(new_n19299), .O(new_n19301));
  nor2 g19108(.a(new_n19301), .b(new_n19268), .O(new_n19302));
  nor2 g19109(.a(new_n19302), .b(new_n19300), .O(new_n19303));
  inv1 g19110(.a(new_n19303), .O(new_n19304));
  nor2 g19111(.a(new_n19304), .b(new_n19258), .O(new_n19305));
  nor2 g19112(.a(new_n19303), .b(new_n19257), .O(new_n19306));
  nor2 g19113(.a(new_n19306), .b(new_n19305), .O(new_n19307));
  inv1 g19114(.a(new_n19307), .O(new_n19308));
  nor2 g19115(.a(new_n19308), .b(new_n19199), .O(new_n19309));
  inv1 g19116(.a(new_n19199), .O(new_n19310));
  nor2 g19117(.a(new_n19307), .b(new_n19310), .O(new_n19311));
  nor2 g19118(.a(new_n19311), .b(new_n19309), .O(new_n19312));
  inv1 g19119(.a(new_n19312), .O(new_n19313));
  nor2 g19120(.a(new_n19313), .b(new_n19198), .O(new_n19314));
  nor2 g19121(.a(new_n19312), .b(new_n19197), .O(new_n19315));
  nor2 g19122(.a(new_n19315), .b(new_n19314), .O(new_n19316));
  inv1 g19123(.a(new_n19316), .O(new_n19317));
  nor2 g19124(.a(new_n19037), .b(new_n18983), .O(new_n19318));
  nor2 g19125(.a(new_n19077), .b(new_n19070), .O(new_n19319));
  inv1 g19126(.a(new_n19319), .O(new_n19320));
  nor2 g19127(.a(new_n19143), .b(new_n19136), .O(new_n19321));
  inv1 g19128(.a(new_n19321), .O(new_n19322));
  nor2 g19129(.a(new_n19322), .b(new_n19320), .O(new_n19323));
  nor2 g19130(.a(new_n19321), .b(new_n19319), .O(new_n19324));
  nor2 g19131(.a(new_n19324), .b(new_n19323), .O(new_n19325));
  nor2 g19132(.a(new_n19134), .b(new_n19126), .O(new_n19326));
  nor2 g19133(.a(new_n19053), .b(new_n19046), .O(new_n19327));
  nor2 g19134(.a(new_n19327), .b(new_n19326), .O(new_n19328));
  inv1 g19135(.a(new_n19326), .O(new_n19329));
  inv1 g19136(.a(new_n19327), .O(new_n19330));
  nor2 g19137(.a(new_n19330), .b(new_n19329), .O(new_n19331));
  nor2 g19138(.a(new_n19331), .b(new_n19328), .O(new_n19332));
  inv1 g19139(.a(new_n19332), .O(new_n19333));
  nor2 g19140(.a(new_n11596), .b(new_n2121), .O(new_n19334));
  inv1 g19141(.a(new_n19334), .O(new_n19335));
  nor2 g19142(.a(new_n6958), .b(new_n4682), .O(new_n19336));
  nor2 g19143(.a(new_n19336), .b(new_n19048), .O(new_n19337));
  nor2 g19144(.a(new_n7294), .b(new_n4682), .O(new_n19338));
  inv1 g19145(.a(new_n19338), .O(new_n19339));
  nor2 g19146(.a(new_n19339), .b(new_n18813), .O(new_n19340));
  nor2 g19147(.a(new_n19340), .b(new_n19337), .O(new_n19341));
  nor2 g19148(.a(new_n19341), .b(new_n19335), .O(new_n19342));
  inv1 g19149(.a(new_n19341), .O(new_n19343));
  nor2 g19150(.a(new_n19343), .b(new_n19334), .O(new_n19344));
  nor2 g19151(.a(new_n19344), .b(new_n19342), .O(new_n19345));
  nor2 g19152(.a(new_n19345), .b(new_n19333), .O(new_n19346));
  inv1 g19153(.a(new_n19345), .O(new_n19347));
  nor2 g19154(.a(new_n19347), .b(new_n19332), .O(new_n19348));
  nor2 g19155(.a(new_n19348), .b(new_n19346), .O(new_n19349));
  nor2 g19156(.a(new_n19349), .b(new_n19325), .O(new_n19350));
  inv1 g19157(.a(new_n19325), .O(new_n19351));
  inv1 g19158(.a(new_n19349), .O(new_n19352));
  nor2 g19159(.a(new_n19352), .b(new_n19351), .O(new_n19353));
  nor2 g19160(.a(new_n19353), .b(new_n19350), .O(new_n19354));
  inv1 g19161(.a(new_n19354), .O(new_n19355));
  nor2 g19162(.a(new_n19146), .b(new_n19094), .O(new_n19356));
  nor2 g19163(.a(new_n19356), .b(new_n19355), .O(new_n19357));
  inv1 g19164(.a(new_n19356), .O(new_n19358));
  nor2 g19165(.a(new_n19358), .b(new_n19354), .O(new_n19359));
  nor2 g19166(.a(new_n19359), .b(new_n19357), .O(new_n19360));
  inv1 g19167(.a(new_n19360), .O(new_n19361));
  nor2 g19168(.a(new_n19361), .b(new_n19318), .O(new_n19362));
  inv1 g19169(.a(new_n19318), .O(new_n19363));
  nor2 g19170(.a(new_n19360), .b(new_n19363), .O(new_n19364));
  nor2 g19171(.a(new_n19364), .b(new_n19362), .O(new_n19365));
  inv1 g19172(.a(new_n19365), .O(new_n19366));
  nor2 g19173(.a(new_n19155), .b(new_n19150), .O(new_n19367));
  nor2 g19174(.a(new_n19367), .b(new_n19366), .O(new_n19368));
  inv1 g19175(.a(new_n19367), .O(new_n19369));
  nor2 g19176(.a(new_n19369), .b(new_n19365), .O(new_n19370));
  nor2 g19177(.a(new_n19370), .b(new_n19368), .O(new_n19371));
  inv1 g19178(.a(new_n19371), .O(new_n19372));
  nor2 g19179(.a(new_n19372), .b(new_n19317), .O(new_n19373));
  nor2 g19180(.a(new_n19371), .b(new_n19316), .O(new_n19374));
  nor2 g19181(.a(new_n19374), .b(new_n19373), .O(new_n19375));
  inv1 g19182(.a(new_n19375), .O(new_n19376));
  nor2 g19183(.a(new_n19161), .b(new_n18976), .O(new_n19377));
  inv1 g19184(.a(new_n19377), .O(new_n19378));
  nor2 g19185(.a(new_n19378), .b(new_n19376), .O(new_n19379));
  nor2 g19186(.a(new_n19377), .b(new_n19375), .O(new_n19380));
  nor2 g19187(.a(new_n19380), .b(new_n19379), .O(new_n19381));
  nor2 g19188(.a(new_n19169), .b(new_n19164), .O(new_n19382));
  nor2 g19189(.a(new_n19382), .b(new_n19165), .O(new_n19383));
  inv1 g19190(.a(new_n19383), .O(new_n19384));
  nor2 g19191(.a(new_n19384), .b(new_n19381), .O(new_n19385));
  inv1 g19192(.a(new_n19381), .O(new_n19386));
  nor2 g19193(.a(new_n19383), .b(new_n19386), .O(new_n19387));
  nor2 g19194(.a(new_n19387), .b(new_n19385), .O(\asquared[90] ));
  nor2 g19195(.a(new_n19373), .b(new_n19368), .O(new_n19389));
  inv1 g19196(.a(new_n19389), .O(new_n19390));
  nor2 g19197(.a(new_n19194), .b(new_n19190), .O(new_n19391));
  inv1 g19198(.a(new_n19391), .O(new_n19392));
  nor2 g19199(.a(new_n19243), .b(new_n5971), .O(new_n19393));
  nor2 g19200(.a(new_n19236), .b(new_n19229), .O(new_n19394));
  nor2 g19201(.a(new_n19394), .b(new_n19393), .O(new_n19395));
  inv1 g19202(.a(new_n19393), .O(new_n19396));
  inv1 g19203(.a(new_n19394), .O(new_n19397));
  nor2 g19204(.a(new_n19397), .b(new_n19396), .O(new_n19398));
  nor2 g19205(.a(new_n19398), .b(new_n19395), .O(new_n19399));
  nor2 g19206(.a(new_n19278), .b(new_n19272), .O(new_n19400));
  nor2 g19207(.a(new_n19400), .b(new_n19399), .O(new_n19401));
  inv1 g19208(.a(new_n19399), .O(new_n19402));
  inv1 g19209(.a(new_n19400), .O(new_n19403));
  nor2 g19210(.a(new_n19403), .b(new_n19402), .O(new_n19404));
  nor2 g19211(.a(new_n19404), .b(new_n19401), .O(new_n19405));
  inv1 g19212(.a(new_n19405), .O(new_n19406));
  nor2 g19213(.a(new_n19251), .b(new_n19245), .O(new_n19407));
  inv1 g19214(.a(new_n19407), .O(new_n19408));
  nor2 g19215(.a(new_n19302), .b(new_n19295), .O(new_n19409));
  inv1 g19216(.a(new_n19409), .O(new_n19410));
  nor2 g19217(.a(new_n19410), .b(new_n19408), .O(new_n19411));
  nor2 g19218(.a(new_n19409), .b(new_n19407), .O(new_n19412));
  nor2 g19219(.a(new_n19412), .b(new_n19411), .O(new_n19413));
  inv1 g19220(.a(new_n19413), .O(new_n19414));
  nor2 g19221(.a(new_n19414), .b(new_n19406), .O(new_n19415));
  nor2 g19222(.a(new_n19413), .b(new_n19405), .O(new_n19416));
  nor2 g19223(.a(new_n19416), .b(new_n19415), .O(new_n19417));
  inv1 g19224(.a(new_n19417), .O(new_n19418));
  nor2 g19225(.a(new_n19305), .b(new_n19255), .O(new_n19419));
  nor2 g19226(.a(new_n19419), .b(new_n19418), .O(new_n19420));
  inv1 g19227(.a(new_n19419), .O(new_n19421));
  nor2 g19228(.a(new_n19421), .b(new_n19417), .O(new_n19422));
  nor2 g19229(.a(new_n19422), .b(new_n19420), .O(new_n19423));
  nor2 g19230(.a(new_n19423), .b(new_n19392), .O(new_n19424));
  inv1 g19231(.a(new_n19423), .O(new_n19425));
  nor2 g19232(.a(new_n19425), .b(new_n19391), .O(new_n19426));
  nor2 g19233(.a(new_n19426), .b(new_n19424), .O(new_n19427));
  nor2 g19234(.a(new_n19314), .b(new_n19309), .O(new_n19428));
  inv1 g19235(.a(new_n19428), .O(new_n19429));
  nor2 g19236(.a(new_n19429), .b(new_n19427), .O(new_n19430));
  inv1 g19237(.a(new_n19427), .O(new_n19431));
  nor2 g19238(.a(new_n19428), .b(new_n19431), .O(new_n19432));
  nor2 g19239(.a(new_n19432), .b(new_n19430), .O(new_n19433));
  nor2 g19240(.a(new_n19362), .b(new_n19357), .O(new_n19434));
  nor2 g19241(.a(new_n19293), .b(new_n19285), .O(new_n19435));
  nor2 g19242(.a(new_n19267), .b(new_n19262), .O(new_n19436));
  nor2 g19243(.a(new_n19436), .b(new_n19435), .O(new_n19437));
  inv1 g19244(.a(new_n19435), .O(new_n19438));
  inv1 g19245(.a(new_n19436), .O(new_n19439));
  nor2 g19246(.a(new_n19439), .b(new_n19438), .O(new_n19440));
  nor2 g19247(.a(new_n19440), .b(new_n19437), .O(new_n19441));
  nor2 g19248(.a(new_n19344), .b(new_n19337), .O(new_n19442));
  nor2 g19249(.a(new_n19442), .b(new_n19441), .O(new_n19443));
  inv1 g19250(.a(new_n19441), .O(new_n19444));
  inv1 g19251(.a(new_n19442), .O(new_n19445));
  nor2 g19252(.a(new_n19445), .b(new_n19444), .O(new_n19446));
  nor2 g19253(.a(new_n19446), .b(new_n19443), .O(new_n19447));
  nor2 g19254(.a(new_n19184), .b(new_n19178), .O(new_n19448));
  inv1 g19255(.a(new_n19448), .O(new_n19449));
  nor2 g19256(.a(new_n19449), .b(new_n19447), .O(new_n19450));
  inv1 g19257(.a(new_n19447), .O(new_n19451));
  nor2 g19258(.a(new_n19448), .b(new_n19451), .O(new_n19452));
  nor2 g19259(.a(new_n19452), .b(new_n19450), .O(new_n19453));
  inv1 g19260(.a(new_n19453), .O(new_n19454));
  nor2 g19261(.a(new_n6893), .b(new_n5178), .O(new_n19455));
  inv1 g19262(.a(new_n19455), .O(new_n19456));
  nor2 g19263(.a(new_n6274), .b(new_n5796), .O(new_n19457));
  nor2 g19264(.a(new_n19457), .b(new_n19230), .O(new_n19458));
  inv1 g19265(.a(new_n19228), .O(new_n19459));
  nor2 g19266(.a(new_n6570), .b(new_n5796), .O(new_n19460));
  inv1 g19267(.a(new_n19460), .O(new_n19461));
  nor2 g19268(.a(new_n19461), .b(new_n19459), .O(new_n19462));
  nor2 g19269(.a(new_n19462), .b(new_n19458), .O(new_n19463));
  nor2 g19270(.a(new_n19463), .b(new_n19456), .O(new_n19464));
  inv1 g19271(.a(new_n19463), .O(new_n19465));
  nor2 g19272(.a(new_n19465), .b(new_n19455), .O(new_n19466));
  nor2 g19273(.a(new_n19466), .b(new_n19464), .O(new_n19467));
  inv1 g19274(.a(new_n19467), .O(new_n19468));
  nor2 g19275(.a(new_n8946), .b(new_n3722), .O(new_n19469));
  nor2 g19276(.a(new_n9658), .b(new_n3231), .O(new_n19470));
  nor2 g19277(.a(new_n9156), .b(new_n3533), .O(new_n19471));
  nor2 g19278(.a(new_n19471), .b(new_n19470), .O(new_n19472));
  nor2 g19279(.a(new_n9658), .b(new_n3533), .O(new_n19473));
  inv1 g19280(.a(new_n19473), .O(new_n19474));
  nor2 g19281(.a(new_n19474), .b(new_n18761), .O(new_n19475));
  nor2 g19282(.a(new_n19475), .b(new_n19472), .O(new_n19476));
  inv1 g19283(.a(new_n19476), .O(new_n19477));
  nor2 g19284(.a(new_n19477), .b(new_n19469), .O(new_n19478));
  inv1 g19285(.a(new_n19469), .O(new_n19479));
  nor2 g19286(.a(new_n19476), .b(new_n19479), .O(new_n19480));
  nor2 g19287(.a(new_n19480), .b(new_n19478), .O(new_n19481));
  nor2 g19288(.a(new_n8476), .b(new_n3870), .O(new_n19482));
  inv1 g19289(.a(new_n19482), .O(new_n19483));
  nor2 g19290(.a(new_n8170), .b(new_n4093), .O(new_n19484));
  nor2 g19291(.a(new_n19484), .b(new_n19287), .O(new_n19485));
  nor2 g19292(.a(new_n8170), .b(new_n4366), .O(new_n19486));
  inv1 g19293(.a(new_n19486), .O(new_n19487));
  nor2 g19294(.a(new_n19487), .b(new_n19104), .O(new_n19488));
  nor2 g19295(.a(new_n19488), .b(new_n19485), .O(new_n19489));
  nor2 g19296(.a(new_n19489), .b(new_n19483), .O(new_n19490));
  inv1 g19297(.a(new_n19489), .O(new_n19491));
  nor2 g19298(.a(new_n19491), .b(new_n19482), .O(new_n19492));
  nor2 g19299(.a(new_n19492), .b(new_n19490), .O(new_n19493));
  nor2 g19300(.a(new_n19493), .b(new_n19481), .O(new_n19494));
  inv1 g19301(.a(new_n19481), .O(new_n19495));
  inv1 g19302(.a(new_n19493), .O(new_n19496));
  nor2 g19303(.a(new_n19496), .b(new_n19495), .O(new_n19497));
  nor2 g19304(.a(new_n19497), .b(new_n19494), .O(new_n19498));
  nor2 g19305(.a(new_n19498), .b(new_n19468), .O(new_n19499));
  inv1 g19306(.a(new_n19498), .O(new_n19500));
  nor2 g19307(.a(new_n19500), .b(new_n19467), .O(new_n19501));
  nor2 g19308(.a(new_n19501), .b(new_n19499), .O(new_n19502));
  inv1 g19309(.a(new_n19502), .O(new_n19503));
  nor2 g19310(.a(new_n19503), .b(new_n19454), .O(new_n19504));
  nor2 g19311(.a(new_n19502), .b(new_n19453), .O(new_n19505));
  nor2 g19312(.a(new_n19505), .b(new_n19504), .O(new_n19506));
  inv1 g19313(.a(new_n19506), .O(new_n19507));
  nor2 g19314(.a(new_n19507), .b(new_n19434), .O(new_n19508));
  inv1 g19315(.a(new_n19434), .O(new_n19509));
  nor2 g19316(.a(new_n19506), .b(new_n19509), .O(new_n19510));
  nor2 g19317(.a(new_n19510), .b(new_n19508), .O(new_n19511));
  inv1 g19318(.a(new_n19511), .O(new_n19512));
  nor2 g19319(.a(new_n19353), .b(new_n19324), .O(new_n19513));
  nor2 g19320(.a(new_n19211), .b(new_n19205), .O(new_n19514));
  nor2 g19321(.a(new_n7537), .b(new_n4425), .O(new_n19515));
  inv1 g19322(.a(new_n19515), .O(new_n19516));
  nor2 g19323(.a(new_n6958), .b(new_n4954), .O(new_n19517));
  nor2 g19324(.a(new_n19517), .b(new_n19338), .O(new_n19518));
  inv1 g19325(.a(new_n19336), .O(new_n19519));
  nor2 g19326(.a(new_n7294), .b(new_n4954), .O(new_n19520));
  inv1 g19327(.a(new_n19520), .O(new_n19521));
  nor2 g19328(.a(new_n19521), .b(new_n19519), .O(new_n19522));
  nor2 g19329(.a(new_n19522), .b(new_n19518), .O(new_n19523));
  nor2 g19330(.a(new_n19523), .b(new_n19516), .O(new_n19524));
  inv1 g19331(.a(new_n19523), .O(new_n19525));
  nor2 g19332(.a(new_n19525), .b(new_n19515), .O(new_n19526));
  nor2 g19333(.a(new_n19526), .b(new_n19524), .O(new_n19527));
  nor2 g19334(.a(new_n19527), .b(new_n19514), .O(new_n19528));
  inv1 g19335(.a(new_n19514), .O(new_n19529));
  inv1 g19336(.a(new_n19527), .O(new_n19530));
  nor2 g19337(.a(new_n19530), .b(new_n19529), .O(new_n19531));
  nor2 g19338(.a(new_n19531), .b(new_n19528), .O(new_n19532));
  nor2 g19339(.a(new_n19346), .b(new_n19331), .O(new_n19533));
  inv1 g19340(.a(new_n19533), .O(new_n19534));
  nor2 g19341(.a(new_n19534), .b(new_n19532), .O(new_n19535));
  inv1 g19342(.a(new_n19532), .O(new_n19536));
  nor2 g19343(.a(new_n19533), .b(new_n19536), .O(new_n19537));
  nor2 g19344(.a(new_n19537), .b(new_n19535), .O(new_n19538));
  inv1 g19345(.a(new_n19538), .O(new_n19539));
  nor2 g19346(.a(new_n11596), .b(new_n2184), .O(new_n19540));
  nor2 g19347(.a(new_n11186), .b(new_n2433), .O(new_n19541));
  nor2 g19348(.a(new_n19541), .b(new_n19217), .O(new_n19542));
  nor2 g19349(.a(new_n11186), .b(new_n2506), .O(new_n19543));
  inv1 g19350(.a(new_n19543), .O(new_n19544));
  nor2 g19351(.a(new_n19544), .b(new_n19117), .O(new_n19545));
  nor2 g19352(.a(new_n19545), .b(new_n19542), .O(new_n19546));
  inv1 g19353(.a(new_n19546), .O(new_n19547));
  nor2 g19354(.a(new_n19547), .b(new_n19540), .O(new_n19548));
  inv1 g19355(.a(new_n19540), .O(new_n19549));
  nor2 g19356(.a(new_n19546), .b(new_n19549), .O(new_n19550));
  nor2 g19357(.a(new_n19550), .b(new_n19548), .O(new_n19551));
  nor2 g19358(.a(new_n19224), .b(new_n19219), .O(new_n19552));
  nor2 g19359(.a(new_n10320), .b(new_n2826), .O(new_n19553));
  nor2 g19360(.a(new_n19553), .b(new_n19062), .O(new_n19554));
  inv1 g19361(.a(new_n19261), .O(new_n19555));
  nor2 g19362(.a(new_n10320), .b(new_n3057), .O(new_n19556));
  inv1 g19363(.a(new_n19556), .O(new_n19557));
  nor2 g19364(.a(new_n19557), .b(new_n19555), .O(new_n19558));
  nor2 g19365(.a(new_n19558), .b(new_n19554), .O(new_n19559));
  nor2 g19366(.a(new_n10468), .b(new_n2660), .O(new_n19560));
  nor2 g19367(.a(new_n19560), .b(new_n19559), .O(new_n19561));
  inv1 g19368(.a(new_n19559), .O(new_n19562));
  inv1 g19369(.a(new_n19560), .O(new_n19563));
  nor2 g19370(.a(new_n19563), .b(new_n19562), .O(new_n19564));
  nor2 g19371(.a(new_n19564), .b(new_n19561), .O(new_n19565));
  inv1 g19372(.a(new_n19565), .O(new_n19566));
  nor2 g19373(.a(new_n19566), .b(new_n19552), .O(new_n19567));
  inv1 g19374(.a(new_n19552), .O(new_n19568));
  nor2 g19375(.a(new_n19565), .b(new_n19568), .O(new_n19569));
  nor2 g19376(.a(new_n19569), .b(new_n19567), .O(new_n19570));
  inv1 g19377(.a(new_n19570), .O(new_n19571));
  nor2 g19378(.a(new_n19571), .b(new_n19551), .O(new_n19572));
  inv1 g19379(.a(new_n19551), .O(new_n19573));
  nor2 g19380(.a(new_n19570), .b(new_n19573), .O(new_n19574));
  nor2 g19381(.a(new_n19574), .b(new_n19572), .O(new_n19575));
  inv1 g19382(.a(new_n19575), .O(new_n19576));
  nor2 g19383(.a(new_n19576), .b(new_n19539), .O(new_n19577));
  nor2 g19384(.a(new_n19575), .b(new_n19538), .O(new_n19578));
  nor2 g19385(.a(new_n19578), .b(new_n19577), .O(new_n19579));
  inv1 g19386(.a(new_n19579), .O(new_n19580));
  nor2 g19387(.a(new_n19580), .b(new_n19513), .O(new_n19581));
  inv1 g19388(.a(new_n19513), .O(new_n19582));
  nor2 g19389(.a(new_n19579), .b(new_n19582), .O(new_n19583));
  nor2 g19390(.a(new_n19583), .b(new_n19581), .O(new_n19584));
  inv1 g19391(.a(new_n19584), .O(new_n19585));
  nor2 g19392(.a(new_n19585), .b(new_n19512), .O(new_n19586));
  nor2 g19393(.a(new_n19584), .b(new_n19511), .O(new_n19587));
  nor2 g19394(.a(new_n19587), .b(new_n19586), .O(new_n19588));
  nor2 g19395(.a(new_n19588), .b(new_n19433), .O(new_n19589));
  inv1 g19396(.a(new_n19433), .O(new_n19590));
  inv1 g19397(.a(new_n19588), .O(new_n19591));
  nor2 g19398(.a(new_n19591), .b(new_n19590), .O(new_n19592));
  nor2 g19399(.a(new_n19592), .b(new_n19589), .O(new_n19593));
  nor2 g19400(.a(new_n19593), .b(new_n19390), .O(new_n19594));
  inv1 g19401(.a(new_n19593), .O(new_n19595));
  nor2 g19402(.a(new_n19595), .b(new_n19389), .O(new_n19596));
  nor2 g19403(.a(new_n19596), .b(new_n19594), .O(new_n19597));
  inv1 g19404(.a(new_n19597), .O(new_n19598));
  nor2 g19405(.a(new_n19384), .b(new_n19379), .O(new_n19599));
  nor2 g19406(.a(new_n19599), .b(new_n19380), .O(new_n19600));
  inv1 g19407(.a(new_n19600), .O(new_n19601));
  nor2 g19408(.a(new_n19601), .b(new_n19598), .O(new_n19602));
  nor2 g19409(.a(new_n19600), .b(new_n19597), .O(new_n19603));
  nor2 g19410(.a(new_n19603), .b(new_n19602), .O(\asquared[91] ));
  nor2 g19411(.a(new_n19592), .b(new_n19432), .O(new_n19605));
  nor2 g19412(.a(new_n19492), .b(new_n19485), .O(new_n19606));
  nor2 g19413(.a(new_n19548), .b(new_n19542), .O(new_n19607));
  nor2 g19414(.a(new_n19607), .b(new_n19606), .O(new_n19608));
  inv1 g19415(.a(new_n19606), .O(new_n19609));
  inv1 g19416(.a(new_n19607), .O(new_n19610));
  nor2 g19417(.a(new_n19610), .b(new_n19609), .O(new_n19611));
  nor2 g19418(.a(new_n19611), .b(new_n19608), .O(new_n19612));
  nor2 g19419(.a(new_n19564), .b(new_n19558), .O(new_n19613));
  inv1 g19420(.a(new_n19613), .O(new_n19614));
  nor2 g19421(.a(new_n19614), .b(new_n19612), .O(new_n19615));
  inv1 g19422(.a(new_n19612), .O(new_n19616));
  nor2 g19423(.a(new_n19613), .b(new_n19616), .O(new_n19617));
  nor2 g19424(.a(new_n19617), .b(new_n19615), .O(new_n19618));
  nor2 g19425(.a(new_n19537), .b(new_n19528), .O(new_n19619));
  inv1 g19426(.a(new_n19619), .O(new_n19620));
  nor2 g19427(.a(new_n19620), .b(new_n19618), .O(new_n19621));
  inv1 g19428(.a(new_n19618), .O(new_n19622));
  nor2 g19429(.a(new_n19619), .b(new_n19622), .O(new_n19623));
  nor2 g19430(.a(new_n19623), .b(new_n19621), .O(new_n19624));
  nor2 g19431(.a(new_n11596), .b(new_n2433), .O(new_n19625));
  nor2 g19432(.a(new_n7537), .b(new_n4682), .O(new_n19626));
  nor2 g19433(.a(new_n19626), .b(new_n19520), .O(new_n19627));
  nor2 g19434(.a(new_n7537), .b(new_n4954), .O(new_n19628));
  inv1 g19435(.a(new_n19628), .O(new_n19629));
  nor2 g19436(.a(new_n19629), .b(new_n19339), .O(new_n19630));
  nor2 g19437(.a(new_n19630), .b(new_n19627), .O(new_n19631));
  inv1 g19438(.a(new_n19631), .O(new_n19632));
  nor2 g19439(.a(new_n19632), .b(new_n19625), .O(new_n19633));
  inv1 g19440(.a(new_n19625), .O(new_n19634));
  nor2 g19441(.a(new_n19631), .b(new_n19634), .O(new_n19635));
  nor2 g19442(.a(new_n19635), .b(new_n19633), .O(new_n19636));
  nor2 g19443(.a(new_n6893), .b(new_n5393), .O(new_n19637));
  nor2 g19444(.a(new_n19637), .b(new_n19460), .O(new_n19638));
  nor2 g19445(.a(new_n6893), .b(new_n5796), .O(new_n19639));
  inv1 g19446(.a(new_n19639), .O(new_n19640));
  nor2 g19447(.a(new_n19640), .b(new_n19231), .O(new_n19641));
  nor2 g19448(.a(new_n19641), .b(new_n19638), .O(new_n19642));
  nor2 g19449(.a(new_n19642), .b(new_n19274), .O(new_n19643));
  inv1 g19450(.a(new_n19642), .O(new_n19644));
  nor2 g19451(.a(new_n19644), .b(new_n19273), .O(new_n19645));
  nor2 g19452(.a(new_n19645), .b(new_n19643), .O(new_n19646));
  nor2 g19453(.a(new_n19646), .b(new_n19636), .O(new_n19647));
  inv1 g19454(.a(new_n19636), .O(new_n19648));
  inv1 g19455(.a(new_n19646), .O(new_n19649));
  nor2 g19456(.a(new_n19649), .b(new_n19648), .O(new_n19650));
  nor2 g19457(.a(new_n19650), .b(new_n19647), .O(new_n19651));
  inv1 g19458(.a(new_n19651), .O(new_n19652));
  nor2 g19459(.a(new_n6274), .b(\a[45] ), .O(new_n19653));
  nor2 g19460(.a(new_n19653), .b(new_n19544), .O(new_n19654));
  inv1 g19461(.a(new_n19653), .O(new_n19655));
  nor2 g19462(.a(new_n19655), .b(new_n19543), .O(new_n19656));
  nor2 g19463(.a(new_n19656), .b(new_n19654), .O(new_n19657));
  nor2 g19464(.a(new_n19657), .b(new_n19652), .O(new_n19658));
  inv1 g19465(.a(new_n19657), .O(new_n19659));
  nor2 g19466(.a(new_n19659), .b(new_n19651), .O(new_n19660));
  nor2 g19467(.a(new_n19660), .b(new_n19658), .O(new_n19661));
  nor2 g19468(.a(new_n19661), .b(new_n19624), .O(new_n19662));
  inv1 g19469(.a(new_n19624), .O(new_n19663));
  inv1 g19470(.a(new_n19661), .O(new_n19664));
  nor2 g19471(.a(new_n19664), .b(new_n19663), .O(new_n19665));
  nor2 g19472(.a(new_n19665), .b(new_n19662), .O(new_n19666));
  inv1 g19473(.a(new_n19666), .O(new_n19667));
  nor2 g19474(.a(new_n19426), .b(new_n19420), .O(new_n19668));
  nor2 g19475(.a(new_n19668), .b(new_n19667), .O(new_n19669));
  inv1 g19476(.a(new_n19668), .O(new_n19670));
  nor2 g19477(.a(new_n19670), .b(new_n19666), .O(new_n19671));
  nor2 g19478(.a(new_n19671), .b(new_n19669), .O(new_n19672));
  inv1 g19479(.a(new_n19672), .O(new_n19673));
  nor2 g19480(.a(new_n19446), .b(new_n19440), .O(new_n19674));
  inv1 g19481(.a(new_n19674), .O(new_n19675));
  nor2 g19482(.a(new_n19404), .b(new_n19398), .O(new_n19676));
  nor2 g19483(.a(new_n6958), .b(new_n5178), .O(new_n19677));
  inv1 g19484(.a(new_n19677), .O(new_n19678));
  nor2 g19485(.a(new_n8946), .b(new_n3870), .O(new_n19679));
  nor2 g19486(.a(new_n19679), .b(new_n19473), .O(new_n19680));
  nor2 g19487(.a(new_n9658), .b(new_n3870), .O(new_n19681));
  inv1 g19488(.a(new_n19681), .O(new_n19682));
  nor2 g19489(.a(new_n19682), .b(new_n19017), .O(new_n19683));
  nor2 g19490(.a(new_n19683), .b(new_n19680), .O(new_n19684));
  nor2 g19491(.a(new_n19684), .b(new_n19678), .O(new_n19685));
  inv1 g19492(.a(new_n19684), .O(new_n19686));
  nor2 g19493(.a(new_n19686), .b(new_n19677), .O(new_n19687));
  nor2 g19494(.a(new_n19687), .b(new_n19685), .O(new_n19688));
  nor2 g19495(.a(new_n19688), .b(new_n19676), .O(new_n19689));
  inv1 g19496(.a(new_n19676), .O(new_n19690));
  inv1 g19497(.a(new_n19688), .O(new_n19691));
  nor2 g19498(.a(new_n19691), .b(new_n19690), .O(new_n19692));
  nor2 g19499(.a(new_n19692), .b(new_n19689), .O(new_n19693));
  nor2 g19500(.a(new_n19693), .b(new_n19675), .O(new_n19694));
  inv1 g19501(.a(new_n19693), .O(new_n19695));
  nor2 g19502(.a(new_n19695), .b(new_n19674), .O(new_n19696));
  nor2 g19503(.a(new_n19696), .b(new_n19694), .O(new_n19697));
  inv1 g19504(.a(new_n19697), .O(new_n19698));
  nor2 g19505(.a(new_n19415), .b(new_n19412), .O(new_n19699));
  nor2 g19506(.a(new_n10468), .b(new_n2826), .O(new_n19700));
  nor2 g19507(.a(new_n9873), .b(new_n3231), .O(new_n19701));
  nor2 g19508(.a(new_n19701), .b(new_n19556), .O(new_n19702));
  nor2 g19509(.a(new_n10320), .b(new_n3231), .O(new_n19703));
  inv1 g19510(.a(new_n19703), .O(new_n19704));
  nor2 g19511(.a(new_n19704), .b(new_n19063), .O(new_n19705));
  nor2 g19512(.a(new_n19705), .b(new_n19702), .O(new_n19706));
  inv1 g19513(.a(new_n19706), .O(new_n19707));
  nor2 g19514(.a(new_n19707), .b(new_n19700), .O(new_n19708));
  inv1 g19515(.a(new_n19700), .O(new_n19709));
  nor2 g19516(.a(new_n19706), .b(new_n19709), .O(new_n19710));
  nor2 g19517(.a(new_n19710), .b(new_n19708), .O(new_n19711));
  inv1 g19518(.a(new_n19711), .O(new_n19712));
  nor2 g19519(.a(new_n8476), .b(new_n4093), .O(new_n19713));
  inv1 g19520(.a(new_n19713), .O(new_n19714));
  nor2 g19521(.a(new_n8026), .b(new_n4425), .O(new_n19715));
  nor2 g19522(.a(new_n19715), .b(new_n19486), .O(new_n19716));
  nor2 g19523(.a(new_n8170), .b(new_n4425), .O(new_n19717));
  inv1 g19524(.a(new_n19717), .O(new_n19718));
  nor2 g19525(.a(new_n19718), .b(new_n19288), .O(new_n19719));
  nor2 g19526(.a(new_n19719), .b(new_n19716), .O(new_n19720));
  nor2 g19527(.a(new_n19720), .b(new_n19714), .O(new_n19721));
  inv1 g19528(.a(new_n19720), .O(new_n19722));
  nor2 g19529(.a(new_n19722), .b(new_n19713), .O(new_n19723));
  nor2 g19530(.a(new_n19723), .b(new_n19721), .O(new_n19724));
  nor2 g19531(.a(new_n19526), .b(new_n19518), .O(new_n19725));
  inv1 g19532(.a(new_n19725), .O(new_n19726));
  nor2 g19533(.a(new_n19726), .b(new_n19724), .O(new_n19727));
  inv1 g19534(.a(new_n19724), .O(new_n19728));
  nor2 g19535(.a(new_n19725), .b(new_n19728), .O(new_n19729));
  nor2 g19536(.a(new_n19729), .b(new_n19727), .O(new_n19730));
  nor2 g19537(.a(new_n19730), .b(new_n19712), .O(new_n19731));
  inv1 g19538(.a(new_n19730), .O(new_n19732));
  nor2 g19539(.a(new_n19732), .b(new_n19711), .O(new_n19733));
  nor2 g19540(.a(new_n19733), .b(new_n19731), .O(new_n19734));
  inv1 g19541(.a(new_n19734), .O(new_n19735));
  nor2 g19542(.a(new_n19735), .b(new_n19699), .O(new_n19736));
  inv1 g19543(.a(new_n19699), .O(new_n19737));
  nor2 g19544(.a(new_n19734), .b(new_n19737), .O(new_n19738));
  nor2 g19545(.a(new_n19738), .b(new_n19736), .O(new_n19739));
  inv1 g19546(.a(new_n19739), .O(new_n19740));
  nor2 g19547(.a(new_n19740), .b(new_n19698), .O(new_n19741));
  nor2 g19548(.a(new_n19739), .b(new_n19697), .O(new_n19742));
  nor2 g19549(.a(new_n19742), .b(new_n19741), .O(new_n19743));
  inv1 g19550(.a(new_n19743), .O(new_n19744));
  nor2 g19551(.a(new_n19744), .b(new_n19673), .O(new_n19745));
  nor2 g19552(.a(new_n19743), .b(new_n19672), .O(new_n19746));
  nor2 g19553(.a(new_n19746), .b(new_n19745), .O(new_n19747));
  inv1 g19554(.a(new_n19747), .O(new_n19748));
  nor2 g19555(.a(new_n19586), .b(new_n19508), .O(new_n19749));
  nor2 g19556(.a(new_n19581), .b(new_n19577), .O(new_n19750));
  nor2 g19557(.a(new_n19504), .b(new_n19452), .O(new_n19751));
  nor2 g19558(.a(new_n10895), .b(new_n2660), .O(new_n19752));
  inv1 g19559(.a(new_n19752), .O(new_n19753));
  nor2 g19560(.a(new_n19466), .b(new_n19458), .O(new_n19754));
  inv1 g19561(.a(new_n19754), .O(new_n19755));
  nor2 g19562(.a(new_n19755), .b(new_n19753), .O(new_n19756));
  nor2 g19563(.a(new_n19754), .b(new_n19752), .O(new_n19757));
  nor2 g19564(.a(new_n19757), .b(new_n19756), .O(new_n19758));
  nor2 g19565(.a(new_n19478), .b(new_n19472), .O(new_n19759));
  nor2 g19566(.a(new_n19759), .b(new_n19758), .O(new_n19760));
  inv1 g19567(.a(new_n19758), .O(new_n19761));
  inv1 g19568(.a(new_n19759), .O(new_n19762));
  nor2 g19569(.a(new_n19762), .b(new_n19761), .O(new_n19763));
  nor2 g19570(.a(new_n19763), .b(new_n19760), .O(new_n19764));
  inv1 g19571(.a(new_n19764), .O(new_n19765));
  nor2 g19572(.a(new_n19572), .b(new_n19567), .O(new_n19766));
  inv1 g19573(.a(new_n19766), .O(new_n19767));
  nor2 g19574(.a(new_n19501), .b(new_n19494), .O(new_n19768));
  inv1 g19575(.a(new_n19768), .O(new_n19769));
  nor2 g19576(.a(new_n19769), .b(new_n19767), .O(new_n19770));
  nor2 g19577(.a(new_n19768), .b(new_n19766), .O(new_n19771));
  nor2 g19578(.a(new_n19771), .b(new_n19770), .O(new_n19772));
  inv1 g19579(.a(new_n19772), .O(new_n19773));
  nor2 g19580(.a(new_n19773), .b(new_n19765), .O(new_n19774));
  nor2 g19581(.a(new_n19772), .b(new_n19764), .O(new_n19775));
  nor2 g19582(.a(new_n19775), .b(new_n19774), .O(new_n19776));
  inv1 g19583(.a(new_n19776), .O(new_n19777));
  nor2 g19584(.a(new_n19777), .b(new_n19751), .O(new_n19778));
  inv1 g19585(.a(new_n19751), .O(new_n19779));
  nor2 g19586(.a(new_n19776), .b(new_n19779), .O(new_n19780));
  nor2 g19587(.a(new_n19780), .b(new_n19778), .O(new_n19781));
  inv1 g19588(.a(new_n19781), .O(new_n19782));
  nor2 g19589(.a(new_n19782), .b(new_n19750), .O(new_n19783));
  inv1 g19590(.a(new_n19750), .O(new_n19784));
  nor2 g19591(.a(new_n19781), .b(new_n19784), .O(new_n19785));
  nor2 g19592(.a(new_n19785), .b(new_n19783), .O(new_n19786));
  inv1 g19593(.a(new_n19786), .O(new_n19787));
  nor2 g19594(.a(new_n19787), .b(new_n19749), .O(new_n19788));
  inv1 g19595(.a(new_n19749), .O(new_n19789));
  nor2 g19596(.a(new_n19786), .b(new_n19789), .O(new_n19790));
  nor2 g19597(.a(new_n19790), .b(new_n19788), .O(new_n19791));
  inv1 g19598(.a(new_n19791), .O(new_n19792));
  nor2 g19599(.a(new_n19792), .b(new_n19748), .O(new_n19793));
  nor2 g19600(.a(new_n19791), .b(new_n19747), .O(new_n19794));
  nor2 g19601(.a(new_n19794), .b(new_n19793), .O(new_n19795));
  inv1 g19602(.a(new_n19795), .O(new_n19796));
  nor2 g19603(.a(new_n19796), .b(new_n19605), .O(new_n19797));
  inv1 g19604(.a(new_n19605), .O(new_n19798));
  nor2 g19605(.a(new_n19795), .b(new_n19798), .O(new_n19799));
  nor2 g19606(.a(new_n19799), .b(new_n19797), .O(new_n19800));
  inv1 g19607(.a(new_n19800), .O(new_n19801));
  nor2 g19608(.a(new_n19602), .b(new_n19596), .O(new_n19802));
  inv1 g19609(.a(new_n19802), .O(new_n19803));
  nor2 g19610(.a(new_n19803), .b(new_n19801), .O(new_n19804));
  nor2 g19611(.a(new_n19802), .b(new_n19800), .O(new_n19805));
  nor2 g19612(.a(new_n19805), .b(new_n19804), .O(new_n19806));
  inv1 g19613(.a(new_n19806), .O(\asquared[92] ));
  nor2 g19614(.a(new_n19783), .b(new_n19778), .O(new_n19808));
  nor2 g19615(.a(new_n19741), .b(new_n19736), .O(new_n19809));
  nor2 g19616(.a(new_n19774), .b(new_n19771), .O(new_n19810));
  nor2 g19617(.a(new_n19763), .b(new_n19756), .O(new_n19811));
  inv1 g19618(.a(new_n19811), .O(new_n19812));
  nor2 g19619(.a(new_n8026), .b(new_n4682), .O(new_n19813));
  nor2 g19620(.a(new_n19813), .b(new_n19628), .O(new_n19814));
  inv1 g19621(.a(new_n19626), .O(new_n19815));
  nor2 g19622(.a(new_n8026), .b(new_n4954), .O(new_n19816));
  inv1 g19623(.a(new_n19816), .O(new_n19817));
  nor2 g19624(.a(new_n19817), .b(new_n19815), .O(new_n19818));
  nor2 g19625(.a(new_n19818), .b(new_n19814), .O(new_n19819));
  nor2 g19626(.a(new_n19819), .b(new_n19718), .O(new_n19820));
  inv1 g19627(.a(new_n19819), .O(new_n19821));
  nor2 g19628(.a(new_n19821), .b(new_n19717), .O(new_n19822));
  nor2 g19629(.a(new_n19822), .b(new_n19820), .O(new_n19823));
  nor2 g19630(.a(new_n10895), .b(new_n2826), .O(new_n19824));
  nor2 g19631(.a(new_n11186), .b(new_n2660), .O(new_n19825));
  nor2 g19632(.a(new_n19825), .b(new_n19824), .O(new_n19826));
  nor2 g19633(.a(new_n11186), .b(new_n2826), .O(new_n19827));
  inv1 g19634(.a(new_n19827), .O(new_n19828));
  nor2 g19635(.a(new_n19828), .b(new_n19753), .O(new_n19829));
  nor2 g19636(.a(new_n19829), .b(new_n19826), .O(new_n19830));
  inv1 g19637(.a(new_n19830), .O(new_n19831));
  nor2 g19638(.a(new_n19656), .b(new_n6274), .O(new_n19832));
  inv1 g19639(.a(new_n19832), .O(new_n19833));
  nor2 g19640(.a(new_n19833), .b(new_n19831), .O(new_n19834));
  nor2 g19641(.a(new_n19832), .b(new_n19830), .O(new_n19835));
  nor2 g19642(.a(new_n19835), .b(new_n19834), .O(new_n19836));
  inv1 g19643(.a(new_n19836), .O(new_n19837));
  nor2 g19644(.a(new_n19837), .b(new_n19823), .O(new_n19838));
  inv1 g19645(.a(new_n19823), .O(new_n19839));
  nor2 g19646(.a(new_n19836), .b(new_n19839), .O(new_n19840));
  nor2 g19647(.a(new_n19840), .b(new_n19838), .O(new_n19841));
  nor2 g19648(.a(new_n19841), .b(new_n19812), .O(new_n19842));
  inv1 g19649(.a(new_n19841), .O(new_n19843));
  nor2 g19650(.a(new_n19843), .b(new_n19811), .O(new_n19844));
  nor2 g19651(.a(new_n19844), .b(new_n19842), .O(new_n19845));
  nor2 g19652(.a(new_n9156), .b(new_n3870), .O(new_n19846));
  inv1 g19653(.a(new_n19846), .O(new_n19847));
  nor2 g19654(.a(new_n19703), .b(new_n16975), .O(new_n19848));
  nor2 g19655(.a(new_n19704), .b(new_n16976), .O(new_n19849));
  nor2 g19656(.a(new_n19849), .b(new_n19848), .O(new_n19850));
  nor2 g19657(.a(new_n19850), .b(new_n19847), .O(new_n19851));
  inv1 g19658(.a(new_n19850), .O(new_n19852));
  nor2 g19659(.a(new_n19852), .b(new_n19846), .O(new_n19853));
  nor2 g19660(.a(new_n19853), .b(new_n19851), .O(new_n19854));
  nor2 g19661(.a(new_n6958), .b(new_n5393), .O(new_n19855));
  inv1 g19662(.a(new_n19855), .O(new_n19856));
  nor2 g19663(.a(new_n6570), .b(new_n5971), .O(new_n19857));
  nor2 g19664(.a(new_n19857), .b(new_n19639), .O(new_n19858));
  nor2 g19665(.a(new_n6893), .b(new_n5971), .O(new_n19859));
  inv1 g19666(.a(new_n19859), .O(new_n19860));
  nor2 g19667(.a(new_n19860), .b(new_n19461), .O(new_n19861));
  nor2 g19668(.a(new_n19861), .b(new_n19858), .O(new_n19862));
  nor2 g19669(.a(new_n19862), .b(new_n19856), .O(new_n19863));
  inv1 g19670(.a(new_n19862), .O(new_n19864));
  nor2 g19671(.a(new_n19864), .b(new_n19855), .O(new_n19865));
  nor2 g19672(.a(new_n19865), .b(new_n19863), .O(new_n19866));
  nor2 g19673(.a(new_n9873), .b(new_n3533), .O(new_n19867));
  inv1 g19674(.a(new_n19867), .O(new_n19868));
  nor2 g19675(.a(new_n7294), .b(new_n5178), .O(new_n19869));
  nor2 g19676(.a(new_n9658), .b(new_n3722), .O(new_n19870));
  nor2 g19677(.a(new_n19870), .b(new_n19869), .O(new_n19871));
  inv1 g19678(.a(new_n19869), .O(new_n19872));
  inv1 g19679(.a(new_n19870), .O(new_n19873));
  nor2 g19680(.a(new_n19873), .b(new_n19872), .O(new_n19874));
  nor2 g19681(.a(new_n19874), .b(new_n19871), .O(new_n19875));
  nor2 g19682(.a(new_n19875), .b(new_n19868), .O(new_n19876));
  inv1 g19683(.a(new_n19875), .O(new_n19877));
  nor2 g19684(.a(new_n19877), .b(new_n19867), .O(new_n19878));
  nor2 g19685(.a(new_n19878), .b(new_n19876), .O(new_n19879));
  nor2 g19686(.a(new_n19879), .b(new_n19866), .O(new_n19880));
  inv1 g19687(.a(new_n19866), .O(new_n19881));
  inv1 g19688(.a(new_n19879), .O(new_n19882));
  nor2 g19689(.a(new_n19882), .b(new_n19881), .O(new_n19883));
  nor2 g19690(.a(new_n19883), .b(new_n19880), .O(new_n19884));
  inv1 g19691(.a(new_n19884), .O(new_n19885));
  nor2 g19692(.a(new_n19885), .b(new_n19854), .O(new_n19886));
  inv1 g19693(.a(new_n19854), .O(new_n19887));
  nor2 g19694(.a(new_n19884), .b(new_n19887), .O(new_n19888));
  nor2 g19695(.a(new_n19888), .b(new_n19886), .O(new_n19889));
  nor2 g19696(.a(new_n19889), .b(new_n19845), .O(new_n19890));
  inv1 g19697(.a(new_n19845), .O(new_n19891));
  inv1 g19698(.a(new_n19889), .O(new_n19892));
  nor2 g19699(.a(new_n19892), .b(new_n19891), .O(new_n19893));
  nor2 g19700(.a(new_n19893), .b(new_n19890), .O(new_n19894));
  inv1 g19701(.a(new_n19894), .O(new_n19895));
  nor2 g19702(.a(new_n19895), .b(new_n19810), .O(new_n19896));
  inv1 g19703(.a(new_n19810), .O(new_n19897));
  nor2 g19704(.a(new_n19894), .b(new_n19897), .O(new_n19898));
  nor2 g19705(.a(new_n19898), .b(new_n19896), .O(new_n19899));
  inv1 g19706(.a(new_n19899), .O(new_n19900));
  nor2 g19707(.a(new_n19900), .b(new_n19809), .O(new_n19901));
  inv1 g19708(.a(new_n19809), .O(new_n19902));
  nor2 g19709(.a(new_n19899), .b(new_n19902), .O(new_n19903));
  nor2 g19710(.a(new_n19903), .b(new_n19901), .O(new_n19904));
  inv1 g19711(.a(new_n19904), .O(new_n19905));
  nor2 g19712(.a(new_n19905), .b(new_n19808), .O(new_n19906));
  inv1 g19713(.a(new_n19808), .O(new_n19907));
  nor2 g19714(.a(new_n19904), .b(new_n19907), .O(new_n19908));
  nor2 g19715(.a(new_n19908), .b(new_n19906), .O(new_n19909));
  inv1 g19716(.a(new_n19909), .O(new_n19910));
  nor2 g19717(.a(new_n19745), .b(new_n19669), .O(new_n19911));
  nor2 g19718(.a(new_n19617), .b(new_n19611), .O(new_n19912));
  inv1 g19719(.a(new_n19912), .O(new_n19913));
  nor2 g19720(.a(new_n19733), .b(new_n19727), .O(new_n19914));
  inv1 g19721(.a(new_n19914), .O(new_n19915));
  nor2 g19722(.a(new_n19915), .b(new_n19913), .O(new_n19916));
  nor2 g19723(.a(new_n19914), .b(new_n19912), .O(new_n19917));
  nor2 g19724(.a(new_n19917), .b(new_n19916), .O(new_n19918));
  nor2 g19725(.a(new_n19658), .b(new_n19647), .O(new_n19919));
  inv1 g19726(.a(new_n19919), .O(new_n19920));
  nor2 g19727(.a(new_n19920), .b(new_n19918), .O(new_n19921));
  inv1 g19728(.a(new_n19918), .O(new_n19922));
  nor2 g19729(.a(new_n19919), .b(new_n19922), .O(new_n19923));
  nor2 g19730(.a(new_n19923), .b(new_n19921), .O(new_n19924));
  inv1 g19731(.a(new_n19924), .O(new_n19925));
  nor2 g19732(.a(new_n19665), .b(new_n19623), .O(new_n19926));
  nor2 g19733(.a(new_n19696), .b(new_n19689), .O(new_n19927));
  nor2 g19734(.a(new_n19723), .b(new_n19716), .O(new_n19928));
  nor2 g19735(.a(new_n19708), .b(new_n19702), .O(new_n19929));
  nor2 g19736(.a(new_n19929), .b(new_n19928), .O(new_n19930));
  inv1 g19737(.a(new_n19928), .O(new_n19931));
  inv1 g19738(.a(new_n19929), .O(new_n19932));
  nor2 g19739(.a(new_n19932), .b(new_n19931), .O(new_n19933));
  nor2 g19740(.a(new_n19933), .b(new_n19930), .O(new_n19934));
  nor2 g19741(.a(new_n19633), .b(new_n19627), .O(new_n19935));
  nor2 g19742(.a(new_n19935), .b(new_n19934), .O(new_n19936));
  inv1 g19743(.a(new_n19934), .O(new_n19937));
  inv1 g19744(.a(new_n19935), .O(new_n19938));
  nor2 g19745(.a(new_n19938), .b(new_n19937), .O(new_n19939));
  nor2 g19746(.a(new_n19939), .b(new_n19936), .O(new_n19940));
  nor2 g19747(.a(new_n19645), .b(new_n19638), .O(new_n19941));
  nor2 g19748(.a(new_n19687), .b(new_n19680), .O(new_n19942));
  nor2 g19749(.a(new_n19942), .b(new_n19941), .O(new_n19943));
  inv1 g19750(.a(new_n19941), .O(new_n19944));
  inv1 g19751(.a(new_n19942), .O(new_n19945));
  nor2 g19752(.a(new_n19945), .b(new_n19944), .O(new_n19946));
  nor2 g19753(.a(new_n19946), .b(new_n19943), .O(new_n19947));
  inv1 g19754(.a(new_n19947), .O(new_n19948));
  nor2 g19755(.a(new_n10468), .b(new_n3057), .O(new_n19949));
  inv1 g19756(.a(new_n19949), .O(new_n19950));
  nor2 g19757(.a(new_n8946), .b(new_n4093), .O(new_n19951));
  nor2 g19758(.a(new_n8476), .b(new_n4366), .O(new_n19952));
  nor2 g19759(.a(new_n19952), .b(new_n19951), .O(new_n19953));
  nor2 g19760(.a(new_n8946), .b(new_n4366), .O(new_n19954));
  inv1 g19761(.a(new_n19954), .O(new_n19955));
  nor2 g19762(.a(new_n19955), .b(new_n19714), .O(new_n19956));
  nor2 g19763(.a(new_n19956), .b(new_n19953), .O(new_n19957));
  nor2 g19764(.a(new_n19957), .b(new_n19950), .O(new_n19958));
  inv1 g19765(.a(new_n19957), .O(new_n19959));
  nor2 g19766(.a(new_n19959), .b(new_n19949), .O(new_n19960));
  nor2 g19767(.a(new_n19960), .b(new_n19958), .O(new_n19961));
  nor2 g19768(.a(new_n19961), .b(new_n19948), .O(new_n19962));
  inv1 g19769(.a(new_n19961), .O(new_n19963));
  nor2 g19770(.a(new_n19963), .b(new_n19947), .O(new_n19964));
  nor2 g19771(.a(new_n19964), .b(new_n19962), .O(new_n19965));
  nor2 g19772(.a(new_n19965), .b(new_n19940), .O(new_n19966));
  inv1 g19773(.a(new_n19940), .O(new_n19967));
  inv1 g19774(.a(new_n19965), .O(new_n19968));
  nor2 g19775(.a(new_n19968), .b(new_n19967), .O(new_n19969));
  nor2 g19776(.a(new_n19969), .b(new_n19966), .O(new_n19970));
  inv1 g19777(.a(new_n19970), .O(new_n19971));
  nor2 g19778(.a(new_n19971), .b(new_n19927), .O(new_n19972));
  inv1 g19779(.a(new_n19927), .O(new_n19973));
  nor2 g19780(.a(new_n19970), .b(new_n19973), .O(new_n19974));
  nor2 g19781(.a(new_n19974), .b(new_n19972), .O(new_n19975));
  inv1 g19782(.a(new_n19975), .O(new_n19976));
  nor2 g19783(.a(new_n19976), .b(new_n19926), .O(new_n19977));
  inv1 g19784(.a(new_n19926), .O(new_n19978));
  nor2 g19785(.a(new_n19975), .b(new_n19978), .O(new_n19979));
  nor2 g19786(.a(new_n19979), .b(new_n19977), .O(new_n19980));
  inv1 g19787(.a(new_n19980), .O(new_n19981));
  nor2 g19788(.a(new_n19981), .b(new_n19925), .O(new_n19982));
  nor2 g19789(.a(new_n19980), .b(new_n19924), .O(new_n19983));
  nor2 g19790(.a(new_n19983), .b(new_n19982), .O(new_n19984));
  inv1 g19791(.a(new_n19984), .O(new_n19985));
  nor2 g19792(.a(new_n19985), .b(new_n19911), .O(new_n19986));
  inv1 g19793(.a(new_n19911), .O(new_n19987));
  nor2 g19794(.a(new_n19984), .b(new_n19987), .O(new_n19988));
  nor2 g19795(.a(new_n19988), .b(new_n19986), .O(new_n19989));
  inv1 g19796(.a(new_n19989), .O(new_n19990));
  nor2 g19797(.a(new_n19990), .b(new_n19910), .O(new_n19991));
  nor2 g19798(.a(new_n19989), .b(new_n19909), .O(new_n19992));
  nor2 g19799(.a(new_n19992), .b(new_n19991), .O(new_n19993));
  nor2 g19800(.a(new_n19793), .b(new_n19788), .O(new_n19994));
  inv1 g19801(.a(new_n19994), .O(new_n19995));
  nor2 g19802(.a(new_n19995), .b(new_n19993), .O(new_n19996));
  inv1 g19803(.a(new_n19993), .O(new_n19997));
  nor2 g19804(.a(new_n19994), .b(new_n19997), .O(new_n19998));
  nor2 g19805(.a(new_n19998), .b(new_n19996), .O(new_n19999));
  inv1 g19806(.a(new_n19999), .O(new_n20000));
  nor2 g19807(.a(new_n19802), .b(new_n19799), .O(new_n20001));
  nor2 g19808(.a(new_n20001), .b(new_n19797), .O(new_n20002));
  nor2 g19809(.a(new_n20002), .b(new_n20000), .O(new_n20003));
  inv1 g19810(.a(new_n20002), .O(new_n20004));
  nor2 g19811(.a(new_n20004), .b(new_n19999), .O(new_n20005));
  nor2 g19812(.a(new_n20005), .b(new_n20003), .O(\asquared[93] ));
  nor2 g19813(.a(new_n19991), .b(new_n19986), .O(new_n20007));
  nor2 g19814(.a(new_n19906), .b(new_n19901), .O(new_n20008));
  inv1 g19815(.a(new_n20008), .O(new_n20009));
  nor2 g19816(.a(new_n19939), .b(new_n19933), .O(new_n20010));
  inv1 g19817(.a(new_n20010), .O(new_n20011));
  nor2 g19818(.a(new_n19962), .b(new_n19946), .O(new_n20012));
  inv1 g19819(.a(new_n20012), .O(new_n20013));
  nor2 g19820(.a(new_n20013), .b(new_n20011), .O(new_n20014));
  nor2 g19821(.a(new_n20012), .b(new_n20010), .O(new_n20015));
  nor2 g19822(.a(new_n20015), .b(new_n20014), .O(new_n20016));
  nor2 g19823(.a(new_n19886), .b(new_n19880), .O(new_n20017));
  inv1 g19824(.a(new_n20017), .O(new_n20018));
  nor2 g19825(.a(new_n20018), .b(new_n20016), .O(new_n20019));
  inv1 g19826(.a(new_n20016), .O(new_n20020));
  nor2 g19827(.a(new_n20017), .b(new_n20020), .O(new_n20021));
  nor2 g19828(.a(new_n20021), .b(new_n20019), .O(new_n20022));
  inv1 g19829(.a(new_n20022), .O(new_n20023));
  nor2 g19830(.a(new_n19972), .b(new_n19969), .O(new_n20024));
  nor2 g19831(.a(new_n20024), .b(new_n20023), .O(new_n20025));
  inv1 g19832(.a(new_n20024), .O(new_n20026));
  nor2 g19833(.a(new_n20026), .b(new_n20022), .O(new_n20027));
  nor2 g19834(.a(new_n20027), .b(new_n20025), .O(new_n20028));
  inv1 g19835(.a(new_n20028), .O(new_n20029));
  nor2 g19836(.a(new_n19844), .b(new_n19838), .O(new_n20030));
  nor2 g19837(.a(new_n19878), .b(new_n19871), .O(new_n20031));
  nor2 g19838(.a(new_n19865), .b(new_n19858), .O(new_n20032));
  nor2 g19839(.a(new_n20032), .b(new_n20031), .O(new_n20033));
  inv1 g19840(.a(new_n20031), .O(new_n20034));
  inv1 g19841(.a(new_n20032), .O(new_n20035));
  nor2 g19842(.a(new_n20035), .b(new_n20034), .O(new_n20036));
  nor2 g19843(.a(new_n20036), .b(new_n20033), .O(new_n20037));
  nor2 g19844(.a(new_n19822), .b(new_n19814), .O(new_n20038));
  nor2 g19845(.a(new_n20038), .b(new_n20037), .O(new_n20039));
  inv1 g19846(.a(new_n20037), .O(new_n20040));
  inv1 g19847(.a(new_n20038), .O(new_n20041));
  nor2 g19848(.a(new_n20041), .b(new_n20040), .O(new_n20042));
  nor2 g19849(.a(new_n20042), .b(new_n20039), .O(new_n20043));
  inv1 g19850(.a(new_n20043), .O(new_n20044));
  nor2 g19851(.a(new_n19853), .b(new_n19848), .O(new_n20045));
  nor2 g19852(.a(new_n19960), .b(new_n19953), .O(new_n20046));
  nor2 g19853(.a(new_n20046), .b(new_n20045), .O(new_n20047));
  inv1 g19854(.a(new_n20045), .O(new_n20048));
  inv1 g19855(.a(new_n20046), .O(new_n20049));
  nor2 g19856(.a(new_n20049), .b(new_n20048), .O(new_n20050));
  nor2 g19857(.a(new_n20050), .b(new_n20047), .O(new_n20051));
  nor2 g19858(.a(new_n19834), .b(new_n19829), .O(new_n20052));
  inv1 g19859(.a(new_n20052), .O(new_n20053));
  nor2 g19860(.a(new_n20053), .b(new_n20051), .O(new_n20054));
  inv1 g19861(.a(new_n20051), .O(new_n20055));
  nor2 g19862(.a(new_n20052), .b(new_n20055), .O(new_n20056));
  nor2 g19863(.a(new_n20056), .b(new_n20054), .O(new_n20057));
  inv1 g19864(.a(new_n20057), .O(new_n20058));
  nor2 g19865(.a(new_n20058), .b(new_n20044), .O(new_n20059));
  nor2 g19866(.a(new_n20057), .b(new_n20043), .O(new_n20060));
  nor2 g19867(.a(new_n20060), .b(new_n20059), .O(new_n20061));
  inv1 g19868(.a(new_n20061), .O(new_n20062));
  nor2 g19869(.a(new_n20062), .b(new_n20030), .O(new_n20063));
  inv1 g19870(.a(new_n20030), .O(new_n20064));
  nor2 g19871(.a(new_n20061), .b(new_n20064), .O(new_n20065));
  nor2 g19872(.a(new_n20065), .b(new_n20063), .O(new_n20066));
  inv1 g19873(.a(new_n20066), .O(new_n20067));
  nor2 g19874(.a(new_n20067), .b(new_n20029), .O(new_n20068));
  nor2 g19875(.a(new_n20066), .b(new_n20028), .O(new_n20069));
  nor2 g19876(.a(new_n20069), .b(new_n20068), .O(new_n20070));
  nor2 g19877(.a(new_n20070), .b(new_n20009), .O(new_n20071));
  inv1 g19878(.a(new_n20070), .O(new_n20072));
  nor2 g19879(.a(new_n20072), .b(new_n20008), .O(new_n20073));
  nor2 g19880(.a(new_n20073), .b(new_n20071), .O(new_n20074));
  inv1 g19881(.a(new_n20074), .O(new_n20075));
  nor2 g19882(.a(new_n19982), .b(new_n19977), .O(new_n20076));
  inv1 g19883(.a(new_n20076), .O(new_n20077));
  nor2 g19884(.a(new_n19896), .b(new_n19893), .O(new_n20078));
  nor2 g19885(.a(new_n19923), .b(new_n19917), .O(new_n20079));
  nor2 g19886(.a(new_n10320), .b(new_n3533), .O(new_n20080));
  inv1 g19887(.a(new_n20080), .O(new_n20081));
  nor2 g19888(.a(new_n8170), .b(new_n4682), .O(new_n20082));
  nor2 g19889(.a(new_n20082), .b(new_n19816), .O(new_n20083));
  inv1 g19890(.a(new_n19813), .O(new_n20084));
  nor2 g19891(.a(new_n8170), .b(new_n4954), .O(new_n20085));
  inv1 g19892(.a(new_n20085), .O(new_n20086));
  nor2 g19893(.a(new_n20086), .b(new_n20084), .O(new_n20087));
  nor2 g19894(.a(new_n20087), .b(new_n20083), .O(new_n20088));
  nor2 g19895(.a(new_n20088), .b(new_n20081), .O(new_n20089));
  inv1 g19896(.a(new_n20088), .O(new_n20090));
  nor2 g19897(.a(new_n20090), .b(new_n20080), .O(new_n20091));
  nor2 g19898(.a(new_n20091), .b(new_n20089), .O(new_n20092));
  nor2 g19899(.a(new_n11596), .b(new_n2660), .O(new_n20093));
  nor2 g19900(.a(new_n10895), .b(new_n3057), .O(new_n20094));
  nor2 g19901(.a(new_n10468), .b(new_n3231), .O(new_n20095));
  nor2 g19902(.a(new_n20095), .b(new_n20094), .O(new_n20096));
  nor2 g19903(.a(new_n10895), .b(new_n3231), .O(new_n20097));
  inv1 g19904(.a(new_n20097), .O(new_n20098));
  nor2 g19905(.a(new_n20098), .b(new_n19950), .O(new_n20099));
  nor2 g19906(.a(new_n20099), .b(new_n20096), .O(new_n20100));
  inv1 g19907(.a(new_n20100), .O(new_n20101));
  nor2 g19908(.a(new_n20101), .b(new_n20093), .O(new_n20102));
  inv1 g19909(.a(new_n20093), .O(new_n20103));
  nor2 g19910(.a(new_n20100), .b(new_n20103), .O(new_n20104));
  nor2 g19911(.a(new_n20104), .b(new_n20102), .O(new_n20105));
  nor2 g19912(.a(new_n9873), .b(new_n3722), .O(new_n20106));
  inv1 g19913(.a(new_n20106), .O(new_n20107));
  nor2 g19914(.a(new_n8476), .b(new_n4425), .O(new_n20108));
  nor2 g19915(.a(new_n20108), .b(new_n19681), .O(new_n20109));
  nor2 g19916(.a(new_n9658), .b(new_n4425), .O(new_n20110));
  inv1 g19917(.a(new_n20110), .O(new_n20111));
  nor2 g19918(.a(new_n20111), .b(new_n19483), .O(new_n20112));
  nor2 g19919(.a(new_n20112), .b(new_n20109), .O(new_n20113));
  nor2 g19920(.a(new_n20113), .b(new_n20107), .O(new_n20114));
  inv1 g19921(.a(new_n20113), .O(new_n20115));
  nor2 g19922(.a(new_n20115), .b(new_n20106), .O(new_n20116));
  nor2 g19923(.a(new_n20116), .b(new_n20114), .O(new_n20117));
  nor2 g19924(.a(new_n20117), .b(new_n20105), .O(new_n20118));
  inv1 g19925(.a(new_n20105), .O(new_n20119));
  inv1 g19926(.a(new_n20117), .O(new_n20120));
  nor2 g19927(.a(new_n20120), .b(new_n20119), .O(new_n20121));
  nor2 g19928(.a(new_n20121), .b(new_n20118), .O(new_n20122));
  inv1 g19929(.a(new_n20122), .O(new_n20123));
  nor2 g19930(.a(new_n20123), .b(new_n20092), .O(new_n20124));
  inv1 g19931(.a(new_n20092), .O(new_n20125));
  nor2 g19932(.a(new_n20122), .b(new_n20125), .O(new_n20126));
  nor2 g19933(.a(new_n20126), .b(new_n20124), .O(new_n20127));
  nor2 g19934(.a(new_n9156), .b(new_n4093), .O(new_n20128));
  nor2 g19935(.a(new_n19954), .b(new_n19859), .O(new_n20129));
  nor2 g19936(.a(new_n8946), .b(new_n5971), .O(new_n20130));
  inv1 g19937(.a(new_n20130), .O(new_n20131));
  nor2 g19938(.a(new_n20131), .b(new_n18351), .O(new_n20132));
  nor2 g19939(.a(new_n20132), .b(new_n20129), .O(new_n20133));
  inv1 g19940(.a(new_n20133), .O(new_n20134));
  nor2 g19941(.a(new_n20134), .b(new_n20128), .O(new_n20135));
  inv1 g19942(.a(new_n20128), .O(new_n20136));
  nor2 g19943(.a(new_n20133), .b(new_n20136), .O(new_n20137));
  nor2 g19944(.a(new_n20137), .b(new_n20135), .O(new_n20138));
  nor2 g19945(.a(new_n7537), .b(new_n5178), .O(new_n20139));
  inv1 g19946(.a(new_n20139), .O(new_n20140));
  nor2 g19947(.a(new_n6958), .b(new_n5796), .O(new_n20141));
  nor2 g19948(.a(new_n7294), .b(new_n5393), .O(new_n20142));
  nor2 g19949(.a(new_n20142), .b(new_n20141), .O(new_n20143));
  nor2 g19950(.a(new_n7294), .b(new_n5796), .O(new_n20144));
  inv1 g19951(.a(new_n20144), .O(new_n20145));
  nor2 g19952(.a(new_n20145), .b(new_n19856), .O(new_n20146));
  nor2 g19953(.a(new_n20146), .b(new_n20143), .O(new_n20147));
  nor2 g19954(.a(new_n20147), .b(new_n20140), .O(new_n20148));
  inv1 g19955(.a(new_n20147), .O(new_n20149));
  nor2 g19956(.a(new_n20149), .b(new_n20139), .O(new_n20150));
  nor2 g19957(.a(new_n20150), .b(new_n20148), .O(new_n20151));
  nor2 g19958(.a(new_n20151), .b(new_n20138), .O(new_n20152));
  inv1 g19959(.a(new_n20138), .O(new_n20153));
  inv1 g19960(.a(new_n20151), .O(new_n20154));
  nor2 g19961(.a(new_n20154), .b(new_n20153), .O(new_n20155));
  nor2 g19962(.a(new_n20155), .b(new_n20152), .O(new_n20156));
  inv1 g19963(.a(new_n20156), .O(new_n20157));
  nor2 g19964(.a(new_n6570), .b(\a[46] ), .O(new_n20158));
  nor2 g19965(.a(new_n20158), .b(new_n19828), .O(new_n20159));
  inv1 g19966(.a(new_n20158), .O(new_n20160));
  nor2 g19967(.a(new_n20160), .b(new_n19827), .O(new_n20161));
  nor2 g19968(.a(new_n20161), .b(new_n20159), .O(new_n20162));
  nor2 g19969(.a(new_n20162), .b(new_n20157), .O(new_n20163));
  inv1 g19970(.a(new_n20162), .O(new_n20164));
  nor2 g19971(.a(new_n20164), .b(new_n20156), .O(new_n20165));
  nor2 g19972(.a(new_n20165), .b(new_n20163), .O(new_n20166));
  nor2 g19973(.a(new_n20166), .b(new_n20127), .O(new_n20167));
  inv1 g19974(.a(new_n20127), .O(new_n20168));
  inv1 g19975(.a(new_n20166), .O(new_n20169));
  nor2 g19976(.a(new_n20169), .b(new_n20168), .O(new_n20170));
  nor2 g19977(.a(new_n20170), .b(new_n20167), .O(new_n20171));
  inv1 g19978(.a(new_n20171), .O(new_n20172));
  nor2 g19979(.a(new_n20172), .b(new_n20079), .O(new_n20173));
  inv1 g19980(.a(new_n20079), .O(new_n20174));
  nor2 g19981(.a(new_n20171), .b(new_n20174), .O(new_n20175));
  nor2 g19982(.a(new_n20175), .b(new_n20173), .O(new_n20176));
  inv1 g19983(.a(new_n20176), .O(new_n20177));
  nor2 g19984(.a(new_n20177), .b(new_n20078), .O(new_n20178));
  inv1 g19985(.a(new_n20078), .O(new_n20179));
  nor2 g19986(.a(new_n20176), .b(new_n20179), .O(new_n20180));
  nor2 g19987(.a(new_n20180), .b(new_n20178), .O(new_n20181));
  nor2 g19988(.a(new_n20181), .b(new_n20077), .O(new_n20182));
  inv1 g19989(.a(new_n20181), .O(new_n20183));
  nor2 g19990(.a(new_n20183), .b(new_n20076), .O(new_n20184));
  nor2 g19991(.a(new_n20184), .b(new_n20182), .O(new_n20185));
  inv1 g19992(.a(new_n20185), .O(new_n20186));
  nor2 g19993(.a(new_n20186), .b(new_n20075), .O(new_n20187));
  nor2 g19994(.a(new_n20185), .b(new_n20074), .O(new_n20188));
  nor2 g19995(.a(new_n20188), .b(new_n20187), .O(new_n20189));
  inv1 g19996(.a(new_n20189), .O(new_n20190));
  nor2 g19997(.a(new_n20190), .b(new_n20007), .O(new_n20191));
  inv1 g19998(.a(new_n20007), .O(new_n20192));
  nor2 g19999(.a(new_n20189), .b(new_n20192), .O(new_n20193));
  nor2 g20000(.a(new_n20193), .b(new_n20191), .O(new_n20194));
  inv1 g20001(.a(new_n20194), .O(new_n20195));
  nor2 g20002(.a(new_n20003), .b(new_n19998), .O(new_n20196));
  inv1 g20003(.a(new_n20196), .O(new_n20197));
  nor2 g20004(.a(new_n20197), .b(new_n20195), .O(new_n20198));
  nor2 g20005(.a(new_n20196), .b(new_n20194), .O(new_n20199));
  nor2 g20006(.a(new_n20199), .b(new_n20198), .O(new_n20200));
  inv1 g20007(.a(new_n20200), .O(\asquared[94] ));
  nor2 g20008(.a(new_n20184), .b(new_n20178), .O(new_n20202));
  inv1 g20009(.a(new_n20202), .O(new_n20203));
  nor2 g20010(.a(new_n20173), .b(new_n20170), .O(new_n20204));
  nor2 g20011(.a(new_n20056), .b(new_n20050), .O(new_n20205));
  inv1 g20012(.a(new_n20205), .O(new_n20206));
  nor2 g20013(.a(new_n20042), .b(new_n20036), .O(new_n20207));
  inv1 g20014(.a(new_n20207), .O(new_n20208));
  nor2 g20015(.a(new_n20208), .b(new_n20206), .O(new_n20209));
  nor2 g20016(.a(new_n20207), .b(new_n20205), .O(new_n20210));
  nor2 g20017(.a(new_n20210), .b(new_n20209), .O(new_n20211));
  nor2 g20018(.a(new_n20124), .b(new_n20118), .O(new_n20212));
  inv1 g20019(.a(new_n20212), .O(new_n20213));
  nor2 g20020(.a(new_n20213), .b(new_n20211), .O(new_n20214));
  inv1 g20021(.a(new_n20211), .O(new_n20215));
  nor2 g20022(.a(new_n20212), .b(new_n20215), .O(new_n20216));
  nor2 g20023(.a(new_n20216), .b(new_n20214), .O(new_n20217));
  inv1 g20024(.a(new_n20217), .O(new_n20218));
  nor2 g20025(.a(new_n20063), .b(new_n20059), .O(new_n20219));
  nor2 g20026(.a(new_n20219), .b(new_n20218), .O(new_n20220));
  inv1 g20027(.a(new_n20219), .O(new_n20221));
  nor2 g20028(.a(new_n20221), .b(new_n20217), .O(new_n20222));
  nor2 g20029(.a(new_n20222), .b(new_n20220), .O(new_n20223));
  inv1 g20030(.a(new_n20223), .O(new_n20224));
  nor2 g20031(.a(new_n20224), .b(new_n20204), .O(new_n20225));
  inv1 g20032(.a(new_n20204), .O(new_n20226));
  nor2 g20033(.a(new_n20223), .b(new_n20226), .O(new_n20227));
  nor2 g20034(.a(new_n20227), .b(new_n20225), .O(new_n20228));
  nor2 g20035(.a(new_n20228), .b(new_n20203), .O(new_n20229));
  inv1 g20036(.a(new_n20228), .O(new_n20230));
  nor2 g20037(.a(new_n20230), .b(new_n20202), .O(new_n20231));
  nor2 g20038(.a(new_n20231), .b(new_n20229), .O(new_n20232));
  nor2 g20039(.a(new_n20068), .b(new_n20025), .O(new_n20233));
  nor2 g20040(.a(new_n20161), .b(new_n6570), .O(new_n20234));
  inv1 g20041(.a(new_n20234), .O(new_n20235));
  nor2 g20042(.a(new_n20235), .b(new_n16293), .O(new_n20236));
  nor2 g20043(.a(new_n20234), .b(new_n16292), .O(new_n20237));
  nor2 g20044(.a(new_n20237), .b(new_n20236), .O(new_n20238));
  nor2 g20045(.a(new_n20135), .b(new_n20129), .O(new_n20239));
  nor2 g20046(.a(new_n20239), .b(new_n20238), .O(new_n20240));
  inv1 g20047(.a(new_n20238), .O(new_n20241));
  inv1 g20048(.a(new_n20239), .O(new_n20242));
  nor2 g20049(.a(new_n20242), .b(new_n20241), .O(new_n20243));
  nor2 g20050(.a(new_n20243), .b(new_n20240), .O(new_n20244));
  nor2 g20051(.a(new_n20163), .b(new_n20152), .O(new_n20245));
  inv1 g20052(.a(new_n20245), .O(new_n20246));
  nor2 g20053(.a(new_n20246), .b(new_n20244), .O(new_n20247));
  inv1 g20054(.a(new_n20244), .O(new_n20248));
  nor2 g20055(.a(new_n20245), .b(new_n20248), .O(new_n20249));
  nor2 g20056(.a(new_n20249), .b(new_n20247), .O(new_n20250));
  inv1 g20057(.a(new_n20250), .O(new_n20251));
  nor2 g20058(.a(new_n20116), .b(new_n20109), .O(new_n20252));
  nor2 g20059(.a(new_n20102), .b(new_n20096), .O(new_n20253));
  nor2 g20060(.a(new_n20253), .b(new_n20252), .O(new_n20254));
  inv1 g20061(.a(new_n20252), .O(new_n20255));
  inv1 g20062(.a(new_n20253), .O(new_n20256));
  nor2 g20063(.a(new_n20256), .b(new_n20255), .O(new_n20257));
  nor2 g20064(.a(new_n20257), .b(new_n20254), .O(new_n20258));
  nor2 g20065(.a(new_n20091), .b(new_n20083), .O(new_n20259));
  nor2 g20066(.a(new_n20259), .b(new_n20258), .O(new_n20260));
  inv1 g20067(.a(new_n20258), .O(new_n20261));
  inv1 g20068(.a(new_n20259), .O(new_n20262));
  nor2 g20069(.a(new_n20262), .b(new_n20261), .O(new_n20263));
  nor2 g20070(.a(new_n20263), .b(new_n20260), .O(new_n20264));
  inv1 g20071(.a(new_n20264), .O(new_n20265));
  nor2 g20072(.a(new_n20265), .b(new_n20251), .O(new_n20266));
  nor2 g20073(.a(new_n20264), .b(new_n20250), .O(new_n20267));
  nor2 g20074(.a(new_n20267), .b(new_n20266), .O(new_n20268));
  inv1 g20075(.a(new_n20268), .O(new_n20269));
  nor2 g20076(.a(new_n20269), .b(new_n20233), .O(new_n20270));
  inv1 g20077(.a(new_n20233), .O(new_n20271));
  nor2 g20078(.a(new_n20268), .b(new_n20271), .O(new_n20272));
  nor2 g20079(.a(new_n20272), .b(new_n20270), .O(new_n20273));
  inv1 g20080(.a(new_n20273), .O(new_n20274));
  nor2 g20081(.a(new_n20021), .b(new_n20015), .O(new_n20275));
  inv1 g20082(.a(new_n20275), .O(new_n20276));
  nor2 g20083(.a(new_n9873), .b(new_n3870), .O(new_n20277));
  nor2 g20084(.a(new_n7537), .b(new_n5393), .O(new_n20278));
  nor2 g20085(.a(new_n20278), .b(new_n20144), .O(new_n20279));
  inv1 g20086(.a(new_n20142), .O(new_n20280));
  nor2 g20087(.a(new_n7537), .b(new_n5796), .O(new_n20281));
  inv1 g20088(.a(new_n20281), .O(new_n20282));
  nor2 g20089(.a(new_n20282), .b(new_n20280), .O(new_n20283));
  nor2 g20090(.a(new_n20283), .b(new_n20279), .O(new_n20284));
  inv1 g20091(.a(new_n20284), .O(new_n20285));
  nor2 g20092(.a(new_n20285), .b(new_n20277), .O(new_n20286));
  inv1 g20093(.a(new_n20277), .O(new_n20287));
  nor2 g20094(.a(new_n20284), .b(new_n20287), .O(new_n20288));
  nor2 g20095(.a(new_n20288), .b(new_n20286), .O(new_n20289));
  nor2 g20096(.a(new_n8476), .b(new_n4682), .O(new_n20290));
  inv1 g20097(.a(new_n20290), .O(new_n20291));
  nor2 g20098(.a(new_n8026), .b(new_n5178), .O(new_n20292));
  nor2 g20099(.a(new_n20292), .b(new_n20085), .O(new_n20293));
  nor2 g20100(.a(new_n8170), .b(new_n5178), .O(new_n20294));
  inv1 g20101(.a(new_n20294), .O(new_n20295));
  nor2 g20102(.a(new_n20295), .b(new_n19817), .O(new_n20296));
  nor2 g20103(.a(new_n20296), .b(new_n20293), .O(new_n20297));
  nor2 g20104(.a(new_n20297), .b(new_n20291), .O(new_n20298));
  inv1 g20105(.a(new_n20297), .O(new_n20299));
  nor2 g20106(.a(new_n20299), .b(new_n20290), .O(new_n20300));
  nor2 g20107(.a(new_n20300), .b(new_n20298), .O(new_n20301));
  nor2 g20108(.a(new_n20301), .b(new_n20289), .O(new_n20302));
  inv1 g20109(.a(new_n20289), .O(new_n20303));
  inv1 g20110(.a(new_n20301), .O(new_n20304));
  nor2 g20111(.a(new_n20304), .b(new_n20303), .O(new_n20305));
  nor2 g20112(.a(new_n20305), .b(new_n20302), .O(new_n20306));
  inv1 g20113(.a(new_n20306), .O(new_n20307));
  nor2 g20114(.a(new_n6958), .b(new_n5971), .O(new_n20308));
  inv1 g20115(.a(new_n20308), .O(new_n20309));
  nor2 g20116(.a(new_n6893), .b(new_n6274), .O(new_n20310));
  nor2 g20117(.a(new_n9156), .b(new_n4366), .O(new_n20311));
  nor2 g20118(.a(new_n20311), .b(new_n20310), .O(new_n20312));
  inv1 g20119(.a(new_n20310), .O(new_n20313));
  inv1 g20120(.a(new_n20311), .O(new_n20314));
  nor2 g20121(.a(new_n20314), .b(new_n20313), .O(new_n20315));
  nor2 g20122(.a(new_n20315), .b(new_n20312), .O(new_n20316));
  nor2 g20123(.a(new_n20316), .b(new_n20309), .O(new_n20317));
  inv1 g20124(.a(new_n20316), .O(new_n20318));
  nor2 g20125(.a(new_n20318), .b(new_n20308), .O(new_n20319));
  nor2 g20126(.a(new_n20319), .b(new_n20317), .O(new_n20320));
  nor2 g20127(.a(new_n20320), .b(new_n20307), .O(new_n20321));
  inv1 g20128(.a(new_n20320), .O(new_n20322));
  nor2 g20129(.a(new_n20322), .b(new_n20306), .O(new_n20323));
  nor2 g20130(.a(new_n20323), .b(new_n20321), .O(new_n20324));
  nor2 g20131(.a(new_n20324), .b(new_n20276), .O(new_n20325));
  inv1 g20132(.a(new_n20324), .O(new_n20326));
  nor2 g20133(.a(new_n20326), .b(new_n20275), .O(new_n20327));
  nor2 g20134(.a(new_n20327), .b(new_n20325), .O(new_n20328));
  inv1 g20135(.a(new_n20328), .O(new_n20329));
  nor2 g20136(.a(new_n9658), .b(new_n4093), .O(new_n20330));
  inv1 g20137(.a(new_n20330), .O(new_n20331));
  nor2 g20138(.a(new_n10468), .b(new_n3533), .O(new_n20332));
  nor2 g20139(.a(new_n8946), .b(new_n4425), .O(new_n20333));
  nor2 g20140(.a(new_n20333), .b(new_n20332), .O(new_n20334));
  inv1 g20141(.a(new_n20332), .O(new_n20335));
  inv1 g20142(.a(new_n20333), .O(new_n20336));
  nor2 g20143(.a(new_n20336), .b(new_n20335), .O(new_n20337));
  nor2 g20144(.a(new_n20337), .b(new_n20334), .O(new_n20338));
  nor2 g20145(.a(new_n20338), .b(new_n20331), .O(new_n20339));
  inv1 g20146(.a(new_n20338), .O(new_n20340));
  nor2 g20147(.a(new_n20340), .b(new_n20330), .O(new_n20341));
  nor2 g20148(.a(new_n20341), .b(new_n20339), .O(new_n20342));
  inv1 g20149(.a(new_n11871), .O(new_n20343));
  nor2 g20150(.a(new_n10320), .b(new_n3722), .O(new_n20344));
  nor2 g20151(.a(new_n20344), .b(new_n20097), .O(new_n20345));
  nor2 g20152(.a(new_n10895), .b(new_n3722), .O(new_n20346));
  inv1 g20153(.a(new_n20346), .O(new_n20347));
  nor2 g20154(.a(new_n20347), .b(new_n19704), .O(new_n20348));
  nor2 g20155(.a(new_n20348), .b(new_n20345), .O(new_n20349));
  nor2 g20156(.a(new_n20349), .b(new_n20343), .O(new_n20350));
  inv1 g20157(.a(new_n20349), .O(new_n20351));
  nor2 g20158(.a(new_n20351), .b(new_n11871), .O(new_n20352));
  nor2 g20159(.a(new_n20352), .b(new_n20350), .O(new_n20353));
  nor2 g20160(.a(new_n20150), .b(new_n20143), .O(new_n20354));
  inv1 g20161(.a(new_n20354), .O(new_n20355));
  nor2 g20162(.a(new_n20355), .b(new_n20353), .O(new_n20356));
  inv1 g20163(.a(new_n20353), .O(new_n20357));
  nor2 g20164(.a(new_n20354), .b(new_n20357), .O(new_n20358));
  nor2 g20165(.a(new_n20358), .b(new_n20356), .O(new_n20359));
  inv1 g20166(.a(new_n20359), .O(new_n20360));
  nor2 g20167(.a(new_n20360), .b(new_n20342), .O(new_n20361));
  inv1 g20168(.a(new_n20342), .O(new_n20362));
  nor2 g20169(.a(new_n20359), .b(new_n20362), .O(new_n20363));
  nor2 g20170(.a(new_n20363), .b(new_n20361), .O(new_n20364));
  inv1 g20171(.a(new_n20364), .O(new_n20365));
  nor2 g20172(.a(new_n20365), .b(new_n20329), .O(new_n20366));
  nor2 g20173(.a(new_n20364), .b(new_n20328), .O(new_n20367));
  nor2 g20174(.a(new_n20367), .b(new_n20366), .O(new_n20368));
  inv1 g20175(.a(new_n20368), .O(new_n20369));
  nor2 g20176(.a(new_n20369), .b(new_n20274), .O(new_n20370));
  nor2 g20177(.a(new_n20368), .b(new_n20273), .O(new_n20371));
  nor2 g20178(.a(new_n20371), .b(new_n20370), .O(new_n20372));
  nor2 g20179(.a(new_n20372), .b(new_n20232), .O(new_n20373));
  inv1 g20180(.a(new_n20232), .O(new_n20374));
  inv1 g20181(.a(new_n20372), .O(new_n20375));
  nor2 g20182(.a(new_n20375), .b(new_n20374), .O(new_n20376));
  nor2 g20183(.a(new_n20376), .b(new_n20373), .O(new_n20377));
  nor2 g20184(.a(new_n20187), .b(new_n20073), .O(new_n20378));
  inv1 g20185(.a(new_n20378), .O(new_n20379));
  nor2 g20186(.a(new_n20379), .b(new_n20377), .O(new_n20380));
  inv1 g20187(.a(new_n20377), .O(new_n20381));
  nor2 g20188(.a(new_n20378), .b(new_n20381), .O(new_n20382));
  nor2 g20189(.a(new_n20382), .b(new_n20380), .O(new_n20383));
  inv1 g20190(.a(new_n20383), .O(new_n20384));
  nor2 g20191(.a(new_n20196), .b(new_n20193), .O(new_n20385));
  nor2 g20192(.a(new_n20385), .b(new_n20191), .O(new_n20386));
  nor2 g20193(.a(new_n20386), .b(new_n20384), .O(new_n20387));
  inv1 g20194(.a(new_n20386), .O(new_n20388));
  nor2 g20195(.a(new_n20388), .b(new_n20383), .O(new_n20389));
  nor2 g20196(.a(new_n20389), .b(new_n20387), .O(\asquared[95] ));
  nor2 g20197(.a(new_n20376), .b(new_n20231), .O(new_n20391));
  nor2 g20198(.a(new_n20370), .b(new_n20270), .O(new_n20392));
  inv1 g20199(.a(new_n20392), .O(new_n20393));
  nor2 g20200(.a(new_n20366), .b(new_n20327), .O(new_n20394));
  nor2 g20201(.a(new_n20243), .b(new_n20236), .O(new_n20395));
  inv1 g20202(.a(new_n20395), .O(new_n20396));
  nor2 g20203(.a(new_n10320), .b(new_n3870), .O(new_n20397));
  nor2 g20204(.a(new_n10468), .b(new_n3722), .O(new_n20398));
  nor2 g20205(.a(new_n20398), .b(new_n20397), .O(new_n20399));
  inv1 g20206(.a(new_n20344), .O(new_n20400));
  nor2 g20207(.a(new_n10468), .b(new_n3870), .O(new_n20401));
  inv1 g20208(.a(new_n20401), .O(new_n20402));
  nor2 g20209(.a(new_n20402), .b(new_n20400), .O(new_n20403));
  nor2 g20210(.a(new_n20403), .b(new_n20399), .O(new_n20404));
  inv1 g20211(.a(new_n20404), .O(new_n20405));
  nor2 g20212(.a(new_n20319), .b(new_n20312), .O(new_n20406));
  inv1 g20213(.a(new_n20406), .O(new_n20407));
  nor2 g20214(.a(new_n20407), .b(new_n20405), .O(new_n20408));
  nor2 g20215(.a(new_n20406), .b(new_n20404), .O(new_n20409));
  nor2 g20216(.a(new_n20409), .b(new_n20408), .O(new_n20410));
  nor2 g20217(.a(new_n20410), .b(new_n20396), .O(new_n20411));
  inv1 g20218(.a(new_n20410), .O(new_n20412));
  nor2 g20219(.a(new_n20412), .b(new_n20395), .O(new_n20413));
  nor2 g20220(.a(new_n20413), .b(new_n20411), .O(new_n20414));
  nor2 g20221(.a(new_n20263), .b(new_n20257), .O(new_n20415));
  inv1 g20222(.a(new_n20415), .O(new_n20416));
  nor2 g20223(.a(new_n20416), .b(new_n20414), .O(new_n20417));
  inv1 g20224(.a(new_n20414), .O(new_n20418));
  nor2 g20225(.a(new_n20415), .b(new_n20418), .O(new_n20419));
  nor2 g20226(.a(new_n20419), .b(new_n20417), .O(new_n20420));
  inv1 g20227(.a(new_n20420), .O(new_n20421));
  nor2 g20228(.a(new_n20266), .b(new_n20249), .O(new_n20422));
  nor2 g20229(.a(new_n20422), .b(new_n20421), .O(new_n20423));
  inv1 g20230(.a(new_n20422), .O(new_n20424));
  nor2 g20231(.a(new_n20424), .b(new_n20420), .O(new_n20425));
  nor2 g20232(.a(new_n20425), .b(new_n20423), .O(new_n20426));
  inv1 g20233(.a(new_n20426), .O(new_n20427));
  nor2 g20234(.a(new_n20427), .b(new_n20394), .O(new_n20428));
  inv1 g20235(.a(new_n20394), .O(new_n20429));
  nor2 g20236(.a(new_n20426), .b(new_n20429), .O(new_n20430));
  nor2 g20237(.a(new_n20430), .b(new_n20428), .O(new_n20431));
  nor2 g20238(.a(new_n20431), .b(new_n20393), .O(new_n20432));
  inv1 g20239(.a(new_n20431), .O(new_n20433));
  nor2 g20240(.a(new_n20433), .b(new_n20392), .O(new_n20434));
  nor2 g20241(.a(new_n20434), .b(new_n20432), .O(new_n20435));
  inv1 g20242(.a(new_n20435), .O(new_n20436));
  nor2 g20243(.a(new_n20225), .b(new_n20220), .O(new_n20437));
  nor2 g20244(.a(new_n20341), .b(new_n20334), .O(new_n20438));
  nor2 g20245(.a(new_n20352), .b(new_n20345), .O(new_n20439));
  nor2 g20246(.a(new_n20439), .b(new_n20438), .O(new_n20440));
  inv1 g20247(.a(new_n20438), .O(new_n20441));
  inv1 g20248(.a(new_n20439), .O(new_n20442));
  nor2 g20249(.a(new_n20442), .b(new_n20441), .O(new_n20443));
  nor2 g20250(.a(new_n20443), .b(new_n20440), .O(new_n20444));
  nor2 g20251(.a(new_n20300), .b(new_n20293), .O(new_n20445));
  nor2 g20252(.a(new_n20445), .b(new_n20444), .O(new_n20446));
  inv1 g20253(.a(new_n20444), .O(new_n20447));
  inv1 g20254(.a(new_n20445), .O(new_n20448));
  nor2 g20255(.a(new_n20448), .b(new_n20447), .O(new_n20449));
  nor2 g20256(.a(new_n20449), .b(new_n20446), .O(new_n20450));
  inv1 g20257(.a(new_n20450), .O(new_n20451));
  nor2 g20258(.a(new_n20321), .b(new_n20302), .O(new_n20452));
  inv1 g20259(.a(new_n20452), .O(new_n20453));
  nor2 g20260(.a(new_n20361), .b(new_n20356), .O(new_n20454));
  inv1 g20261(.a(new_n20454), .O(new_n20455));
  nor2 g20262(.a(new_n20455), .b(new_n20453), .O(new_n20456));
  nor2 g20263(.a(new_n20454), .b(new_n20452), .O(new_n20457));
  nor2 g20264(.a(new_n20457), .b(new_n20456), .O(new_n20458));
  inv1 g20265(.a(new_n20458), .O(new_n20459));
  nor2 g20266(.a(new_n20459), .b(new_n20451), .O(new_n20460));
  nor2 g20267(.a(new_n20458), .b(new_n20450), .O(new_n20461));
  nor2 g20268(.a(new_n20461), .b(new_n20460), .O(new_n20462));
  inv1 g20269(.a(new_n20462), .O(new_n20463));
  nor2 g20270(.a(new_n20463), .b(new_n20437), .O(new_n20464));
  inv1 g20271(.a(new_n20437), .O(new_n20465));
  nor2 g20272(.a(new_n20462), .b(new_n20465), .O(new_n20466));
  nor2 g20273(.a(new_n20466), .b(new_n20464), .O(new_n20467));
  inv1 g20274(.a(new_n20467), .O(new_n20468));
  nor2 g20275(.a(new_n20216), .b(new_n20210), .O(new_n20469));
  inv1 g20276(.a(new_n20469), .O(new_n20470));
  nor2 g20277(.a(new_n8026), .b(new_n5393), .O(new_n20471));
  nor2 g20278(.a(new_n20471), .b(new_n20281), .O(new_n20472));
  inv1 g20279(.a(new_n20278), .O(new_n20473));
  nor2 g20280(.a(new_n8026), .b(new_n5796), .O(new_n20474));
  inv1 g20281(.a(new_n20474), .O(new_n20475));
  nor2 g20282(.a(new_n20475), .b(new_n20473), .O(new_n20476));
  nor2 g20283(.a(new_n20476), .b(new_n20472), .O(new_n20477));
  nor2 g20284(.a(new_n20477), .b(new_n20295), .O(new_n20478));
  inv1 g20285(.a(new_n20477), .O(new_n20479));
  nor2 g20286(.a(new_n20479), .b(new_n20294), .O(new_n20480));
  nor2 g20287(.a(new_n20480), .b(new_n20478), .O(new_n20481));
  inv1 g20288(.a(new_n20481), .O(new_n20482));
  nor2 g20289(.a(new_n9156), .b(new_n4425), .O(new_n20483));
  inv1 g20290(.a(new_n20483), .O(new_n20484));
  nor2 g20291(.a(new_n6958), .b(new_n6274), .O(new_n20485));
  nor2 g20292(.a(new_n7294), .b(new_n5971), .O(new_n20486));
  nor2 g20293(.a(new_n20486), .b(new_n20485), .O(new_n20487));
  nor2 g20294(.a(new_n7294), .b(new_n6274), .O(new_n20488));
  inv1 g20295(.a(new_n20488), .O(new_n20489));
  nor2 g20296(.a(new_n20489), .b(new_n20309), .O(new_n20490));
  nor2 g20297(.a(new_n20490), .b(new_n20487), .O(new_n20491));
  nor2 g20298(.a(new_n20491), .b(new_n20484), .O(new_n20492));
  inv1 g20299(.a(new_n20491), .O(new_n20493));
  nor2 g20300(.a(new_n20493), .b(new_n20483), .O(new_n20494));
  nor2 g20301(.a(new_n20494), .b(new_n20492), .O(new_n20495));
  nor2 g20302(.a(new_n11186), .b(new_n3231), .O(new_n20496));
  inv1 g20303(.a(new_n20496), .O(new_n20497));
  nor2 g20304(.a(new_n6893), .b(\a[47] ), .O(new_n20498));
  nor2 g20305(.a(new_n20498), .b(new_n20497), .O(new_n20499));
  inv1 g20306(.a(new_n20498), .O(new_n20500));
  nor2 g20307(.a(new_n20500), .b(new_n20496), .O(new_n20501));
  nor2 g20308(.a(new_n20501), .b(new_n20499), .O(new_n20502));
  nor2 g20309(.a(new_n20502), .b(new_n20495), .O(new_n20503));
  inv1 g20310(.a(new_n20495), .O(new_n20504));
  inv1 g20311(.a(new_n20502), .O(new_n20505));
  nor2 g20312(.a(new_n20505), .b(new_n20504), .O(new_n20506));
  nor2 g20313(.a(new_n20506), .b(new_n20503), .O(new_n20507));
  nor2 g20314(.a(new_n20507), .b(new_n20482), .O(new_n20508));
  inv1 g20315(.a(new_n20507), .O(new_n20509));
  nor2 g20316(.a(new_n20509), .b(new_n20481), .O(new_n20510));
  nor2 g20317(.a(new_n20510), .b(new_n20508), .O(new_n20511));
  nor2 g20318(.a(new_n20511), .b(new_n20470), .O(new_n20512));
  inv1 g20319(.a(new_n20511), .O(new_n20513));
  nor2 g20320(.a(new_n20513), .b(new_n20469), .O(new_n20514));
  nor2 g20321(.a(new_n20514), .b(new_n20512), .O(new_n20515));
  inv1 g20322(.a(new_n20515), .O(new_n20516));
  nor2 g20323(.a(new_n8476), .b(new_n4954), .O(new_n20517));
  nor2 g20324(.a(new_n11596), .b(new_n3057), .O(new_n20518));
  nor2 g20325(.a(new_n10895), .b(new_n3533), .O(new_n20519));
  nor2 g20326(.a(new_n20519), .b(new_n20518), .O(new_n20520));
  inv1 g20327(.a(new_n20094), .O(new_n20521));
  nor2 g20328(.a(new_n11596), .b(new_n3533), .O(new_n20522));
  inv1 g20329(.a(new_n20522), .O(new_n20523));
  nor2 g20330(.a(new_n20523), .b(new_n20521), .O(new_n20524));
  nor2 g20331(.a(new_n20524), .b(new_n20520), .O(new_n20525));
  inv1 g20332(.a(new_n20525), .O(new_n20526));
  nor2 g20333(.a(new_n20526), .b(new_n20517), .O(new_n20527));
  inv1 g20334(.a(new_n20517), .O(new_n20528));
  nor2 g20335(.a(new_n20525), .b(new_n20528), .O(new_n20529));
  nor2 g20336(.a(new_n20529), .b(new_n20527), .O(new_n20530));
  inv1 g20337(.a(new_n20530), .O(new_n20531));
  nor2 g20338(.a(new_n9873), .b(new_n4093), .O(new_n20532));
  inv1 g20339(.a(new_n20532), .O(new_n20533));
  nor2 g20340(.a(new_n9658), .b(new_n4366), .O(new_n20534));
  nor2 g20341(.a(new_n8946), .b(new_n4682), .O(new_n20535));
  nor2 g20342(.a(new_n20535), .b(new_n20534), .O(new_n20536));
  nor2 g20343(.a(new_n9658), .b(new_n4682), .O(new_n20537));
  inv1 g20344(.a(new_n20537), .O(new_n20538));
  nor2 g20345(.a(new_n20538), .b(new_n19955), .O(new_n20539));
  nor2 g20346(.a(new_n20539), .b(new_n20536), .O(new_n20540));
  nor2 g20347(.a(new_n20540), .b(new_n20533), .O(new_n20541));
  inv1 g20348(.a(new_n20540), .O(new_n20542));
  nor2 g20349(.a(new_n20542), .b(new_n20532), .O(new_n20543));
  nor2 g20350(.a(new_n20543), .b(new_n20541), .O(new_n20544));
  nor2 g20351(.a(new_n20286), .b(new_n20279), .O(new_n20545));
  inv1 g20352(.a(new_n20545), .O(new_n20546));
  nor2 g20353(.a(new_n20546), .b(new_n20544), .O(new_n20547));
  inv1 g20354(.a(new_n20544), .O(new_n20548));
  nor2 g20355(.a(new_n20545), .b(new_n20548), .O(new_n20549));
  nor2 g20356(.a(new_n20549), .b(new_n20547), .O(new_n20550));
  nor2 g20357(.a(new_n20550), .b(new_n20531), .O(new_n20551));
  inv1 g20358(.a(new_n20550), .O(new_n20552));
  nor2 g20359(.a(new_n20552), .b(new_n20530), .O(new_n20553));
  nor2 g20360(.a(new_n20553), .b(new_n20551), .O(new_n20554));
  inv1 g20361(.a(new_n20554), .O(new_n20555));
  nor2 g20362(.a(new_n20555), .b(new_n20516), .O(new_n20556));
  nor2 g20363(.a(new_n20554), .b(new_n20515), .O(new_n20557));
  nor2 g20364(.a(new_n20557), .b(new_n20556), .O(new_n20558));
  inv1 g20365(.a(new_n20558), .O(new_n20559));
  nor2 g20366(.a(new_n20559), .b(new_n20468), .O(new_n20560));
  nor2 g20367(.a(new_n20558), .b(new_n20467), .O(new_n20561));
  nor2 g20368(.a(new_n20561), .b(new_n20560), .O(new_n20562));
  inv1 g20369(.a(new_n20562), .O(new_n20563));
  nor2 g20370(.a(new_n20563), .b(new_n20436), .O(new_n20564));
  nor2 g20371(.a(new_n20562), .b(new_n20435), .O(new_n20565));
  nor2 g20372(.a(new_n20565), .b(new_n20564), .O(new_n20566));
  inv1 g20373(.a(new_n20566), .O(new_n20567));
  nor2 g20374(.a(new_n20567), .b(new_n20391), .O(new_n20568));
  inv1 g20375(.a(new_n20391), .O(new_n20569));
  nor2 g20376(.a(new_n20566), .b(new_n20569), .O(new_n20570));
  nor2 g20377(.a(new_n20570), .b(new_n20568), .O(new_n20571));
  inv1 g20378(.a(new_n20571), .O(new_n20572));
  nor2 g20379(.a(new_n20387), .b(new_n20382), .O(new_n20573));
  nor2 g20380(.a(new_n20573), .b(new_n20572), .O(new_n20574));
  inv1 g20381(.a(new_n20573), .O(new_n20575));
  nor2 g20382(.a(new_n20575), .b(new_n20571), .O(new_n20576));
  nor2 g20383(.a(new_n20576), .b(new_n20574), .O(\asquared[96] ));
  nor2 g20384(.a(new_n20428), .b(new_n20423), .O(new_n20578));
  nor2 g20385(.a(new_n20501), .b(new_n6893), .O(new_n20579));
  nor2 g20386(.a(new_n20494), .b(new_n20487), .O(new_n20580));
  nor2 g20387(.a(new_n20580), .b(new_n20579), .O(new_n20581));
  inv1 g20388(.a(new_n20579), .O(new_n20582));
  inv1 g20389(.a(new_n20580), .O(new_n20583));
  nor2 g20390(.a(new_n20583), .b(new_n20582), .O(new_n20584));
  nor2 g20391(.a(new_n20584), .b(new_n20581), .O(new_n20585));
  nor2 g20392(.a(new_n20480), .b(new_n20472), .O(new_n20586));
  nor2 g20393(.a(new_n20586), .b(new_n20585), .O(new_n20587));
  inv1 g20394(.a(new_n20585), .O(new_n20588));
  inv1 g20395(.a(new_n20586), .O(new_n20589));
  nor2 g20396(.a(new_n20589), .b(new_n20588), .O(new_n20590));
  nor2 g20397(.a(new_n20590), .b(new_n20587), .O(new_n20591));
  inv1 g20398(.a(new_n20591), .O(new_n20592));
  nor2 g20399(.a(new_n20510), .b(new_n20503), .O(new_n20593));
  inv1 g20400(.a(new_n20593), .O(new_n20594));
  nor2 g20401(.a(new_n20553), .b(new_n20547), .O(new_n20595));
  inv1 g20402(.a(new_n20595), .O(new_n20596));
  nor2 g20403(.a(new_n20596), .b(new_n20594), .O(new_n20597));
  nor2 g20404(.a(new_n20595), .b(new_n20593), .O(new_n20598));
  nor2 g20405(.a(new_n20598), .b(new_n20597), .O(new_n20599));
  inv1 g20406(.a(new_n20599), .O(new_n20600));
  nor2 g20407(.a(new_n20600), .b(new_n20592), .O(new_n20601));
  nor2 g20408(.a(new_n20599), .b(new_n20591), .O(new_n20602));
  nor2 g20409(.a(new_n20602), .b(new_n20601), .O(new_n20603));
  inv1 g20410(.a(new_n20603), .O(new_n20604));
  nor2 g20411(.a(new_n20604), .b(new_n20578), .O(new_n20605));
  inv1 g20412(.a(new_n20578), .O(new_n20606));
  nor2 g20413(.a(new_n20603), .b(new_n20606), .O(new_n20607));
  nor2 g20414(.a(new_n20607), .b(new_n20605), .O(new_n20608));
  inv1 g20415(.a(new_n20608), .O(new_n20609));
  nor2 g20416(.a(new_n20449), .b(new_n20443), .O(new_n20610));
  inv1 g20417(.a(new_n20610), .O(new_n20611));
  nor2 g20418(.a(new_n11596), .b(new_n3231), .O(new_n20612));
  nor2 g20419(.a(new_n11186), .b(new_n3533), .O(new_n20613));
  nor2 g20420(.a(new_n20613), .b(new_n20346), .O(new_n20614));
  inv1 g20421(.a(new_n20519), .O(new_n20615));
  nor2 g20422(.a(new_n11186), .b(new_n3722), .O(new_n20616));
  inv1 g20423(.a(new_n20616), .O(new_n20617));
  nor2 g20424(.a(new_n20617), .b(new_n20615), .O(new_n20618));
  nor2 g20425(.a(new_n20618), .b(new_n20614), .O(new_n20619));
  inv1 g20426(.a(new_n20619), .O(new_n20620));
  nor2 g20427(.a(new_n20620), .b(new_n20612), .O(new_n20621));
  inv1 g20428(.a(new_n20612), .O(new_n20622));
  nor2 g20429(.a(new_n20619), .b(new_n20622), .O(new_n20623));
  nor2 g20430(.a(new_n20623), .b(new_n20621), .O(new_n20624));
  nor2 g20431(.a(new_n8946), .b(new_n4954), .O(new_n20625));
  inv1 g20432(.a(new_n20625), .O(new_n20626));
  nor2 g20433(.a(new_n8476), .b(new_n5178), .O(new_n20627));
  nor2 g20434(.a(new_n8170), .b(new_n5393), .O(new_n20628));
  nor2 g20435(.a(new_n20628), .b(new_n20627), .O(new_n20629));
  nor2 g20436(.a(new_n8476), .b(new_n5393), .O(new_n20630));
  inv1 g20437(.a(new_n20630), .O(new_n20631));
  nor2 g20438(.a(new_n20631), .b(new_n20295), .O(new_n20632));
  nor2 g20439(.a(new_n20632), .b(new_n20629), .O(new_n20633));
  nor2 g20440(.a(new_n20633), .b(new_n20626), .O(new_n20634));
  inv1 g20441(.a(new_n20633), .O(new_n20635));
  nor2 g20442(.a(new_n20635), .b(new_n20625), .O(new_n20636));
  nor2 g20443(.a(new_n20636), .b(new_n20634), .O(new_n20637));
  nor2 g20444(.a(new_n20637), .b(new_n20624), .O(new_n20638));
  inv1 g20445(.a(new_n20624), .O(new_n20639));
  inv1 g20446(.a(new_n20637), .O(new_n20640));
  nor2 g20447(.a(new_n20640), .b(new_n20639), .O(new_n20641));
  nor2 g20448(.a(new_n20641), .b(new_n20638), .O(new_n20642));
  nor2 g20449(.a(new_n20642), .b(new_n20611), .O(new_n20643));
  inv1 g20450(.a(new_n20642), .O(new_n20644));
  nor2 g20451(.a(new_n20644), .b(new_n20610), .O(new_n20645));
  nor2 g20452(.a(new_n20645), .b(new_n20643), .O(new_n20646));
  inv1 g20453(.a(new_n20646), .O(new_n20647));
  nor2 g20454(.a(new_n20543), .b(new_n20536), .O(new_n20648));
  nor2 g20455(.a(new_n20527), .b(new_n20520), .O(new_n20649));
  nor2 g20456(.a(new_n20649), .b(new_n20648), .O(new_n20650));
  inv1 g20457(.a(new_n20648), .O(new_n20651));
  inv1 g20458(.a(new_n20649), .O(new_n20652));
  nor2 g20459(.a(new_n20652), .b(new_n20651), .O(new_n20653));
  nor2 g20460(.a(new_n20653), .b(new_n20650), .O(new_n20654));
  nor2 g20461(.a(new_n20408), .b(new_n20403), .O(new_n20655));
  inv1 g20462(.a(new_n20655), .O(new_n20656));
  nor2 g20463(.a(new_n20656), .b(new_n20654), .O(new_n20657));
  inv1 g20464(.a(new_n20654), .O(new_n20658));
  nor2 g20465(.a(new_n20655), .b(new_n20658), .O(new_n20659));
  nor2 g20466(.a(new_n20659), .b(new_n20657), .O(new_n20660));
  nor2 g20467(.a(new_n20419), .b(new_n20413), .O(new_n20661));
  inv1 g20468(.a(new_n20661), .O(new_n20662));
  nor2 g20469(.a(new_n20662), .b(new_n20660), .O(new_n20663));
  inv1 g20470(.a(new_n20660), .O(new_n20664));
  nor2 g20471(.a(new_n20661), .b(new_n20664), .O(new_n20665));
  nor2 g20472(.a(new_n20665), .b(new_n20663), .O(new_n20666));
  inv1 g20473(.a(new_n20666), .O(new_n20667));
  nor2 g20474(.a(new_n20667), .b(new_n20647), .O(new_n20668));
  nor2 g20475(.a(new_n20666), .b(new_n20646), .O(new_n20669));
  nor2 g20476(.a(new_n20669), .b(new_n20668), .O(new_n20670));
  inv1 g20477(.a(new_n20670), .O(new_n20671));
  nor2 g20478(.a(new_n20671), .b(new_n20609), .O(new_n20672));
  nor2 g20479(.a(new_n20670), .b(new_n20608), .O(new_n20673));
  nor2 g20480(.a(new_n20673), .b(new_n20672), .O(new_n20674));
  inv1 g20481(.a(new_n20674), .O(new_n20675));
  nor2 g20482(.a(new_n20460), .b(new_n20457), .O(new_n20676));
  nor2 g20483(.a(new_n10320), .b(new_n4093), .O(new_n20677));
  nor2 g20484(.a(new_n9156), .b(new_n4682), .O(new_n20678));
  nor2 g20485(.a(new_n20678), .b(new_n20677), .O(new_n20679));
  nor2 g20486(.a(new_n10320), .b(new_n4682), .O(new_n20680));
  inv1 g20487(.a(new_n20680), .O(new_n20681));
  nor2 g20488(.a(new_n20681), .b(new_n20136), .O(new_n20682));
  nor2 g20489(.a(new_n20682), .b(new_n20679), .O(new_n20683));
  inv1 g20490(.a(new_n20683), .O(new_n20684));
  nor2 g20491(.a(new_n20684), .b(new_n20401), .O(new_n20685));
  nor2 g20492(.a(new_n20683), .b(new_n20402), .O(new_n20686));
  nor2 g20493(.a(new_n20686), .b(new_n20685), .O(new_n20687));
  nor2 g20494(.a(new_n9873), .b(new_n4366), .O(new_n20688));
  nor2 g20495(.a(new_n20688), .b(new_n20110), .O(new_n20689));
  inv1 g20496(.a(new_n20534), .O(new_n20690));
  nor2 g20497(.a(new_n9873), .b(new_n4425), .O(new_n20691));
  inv1 g20498(.a(new_n20691), .O(new_n20692));
  nor2 g20499(.a(new_n20692), .b(new_n20690), .O(new_n20693));
  nor2 g20500(.a(new_n20693), .b(new_n20689), .O(new_n20694));
  nor2 g20501(.a(new_n20694), .b(new_n20475), .O(new_n20695));
  inv1 g20502(.a(new_n20694), .O(new_n20696));
  nor2 g20503(.a(new_n20696), .b(new_n20474), .O(new_n20697));
  nor2 g20504(.a(new_n20697), .b(new_n20695), .O(new_n20698));
  nor2 g20505(.a(new_n20698), .b(new_n20687), .O(new_n20699));
  inv1 g20506(.a(new_n20687), .O(new_n20700));
  inv1 g20507(.a(new_n20698), .O(new_n20701));
  nor2 g20508(.a(new_n20701), .b(new_n20700), .O(new_n20702));
  nor2 g20509(.a(new_n20702), .b(new_n20699), .O(new_n20703));
  inv1 g20510(.a(new_n20703), .O(new_n20704));
  nor2 g20511(.a(new_n7537), .b(new_n5971), .O(new_n20705));
  inv1 g20512(.a(new_n20705), .O(new_n20706));
  nor2 g20513(.a(new_n6958), .b(new_n6570), .O(new_n20707));
  nor2 g20514(.a(new_n20707), .b(new_n20488), .O(new_n20708));
  inv1 g20515(.a(new_n20485), .O(new_n20709));
  nor2 g20516(.a(new_n7294), .b(new_n6570), .O(new_n20710));
  inv1 g20517(.a(new_n20710), .O(new_n20711));
  nor2 g20518(.a(new_n20711), .b(new_n20709), .O(new_n20712));
  nor2 g20519(.a(new_n20712), .b(new_n20708), .O(new_n20713));
  nor2 g20520(.a(new_n20713), .b(new_n20706), .O(new_n20714));
  inv1 g20521(.a(new_n20713), .O(new_n20715));
  nor2 g20522(.a(new_n20715), .b(new_n20705), .O(new_n20716));
  nor2 g20523(.a(new_n20716), .b(new_n20714), .O(new_n20717));
  nor2 g20524(.a(new_n20717), .b(new_n20704), .O(new_n20718));
  inv1 g20525(.a(new_n20717), .O(new_n20719));
  nor2 g20526(.a(new_n20719), .b(new_n20703), .O(new_n20720));
  nor2 g20527(.a(new_n20720), .b(new_n20718), .O(new_n20721));
  inv1 g20528(.a(new_n20721), .O(new_n20722));
  nor2 g20529(.a(new_n20722), .b(new_n20676), .O(new_n20723));
  inv1 g20530(.a(new_n20676), .O(new_n20724));
  nor2 g20531(.a(new_n20721), .b(new_n20724), .O(new_n20725));
  nor2 g20532(.a(new_n20725), .b(new_n20723), .O(new_n20726));
  inv1 g20533(.a(new_n20726), .O(new_n20727));
  nor2 g20534(.a(new_n20556), .b(new_n20514), .O(new_n20728));
  nor2 g20535(.a(new_n20728), .b(new_n20727), .O(new_n20729));
  inv1 g20536(.a(new_n20728), .O(new_n20730));
  nor2 g20537(.a(new_n20730), .b(new_n20726), .O(new_n20731));
  nor2 g20538(.a(new_n20731), .b(new_n20729), .O(new_n20732));
  inv1 g20539(.a(new_n20732), .O(new_n20733));
  nor2 g20540(.a(new_n20560), .b(new_n20464), .O(new_n20734));
  nor2 g20541(.a(new_n20734), .b(new_n20733), .O(new_n20735));
  inv1 g20542(.a(new_n20734), .O(new_n20736));
  nor2 g20543(.a(new_n20736), .b(new_n20732), .O(new_n20737));
  nor2 g20544(.a(new_n20737), .b(new_n20735), .O(new_n20738));
  inv1 g20545(.a(new_n20738), .O(new_n20739));
  nor2 g20546(.a(new_n20739), .b(new_n20675), .O(new_n20740));
  nor2 g20547(.a(new_n20738), .b(new_n20674), .O(new_n20741));
  nor2 g20548(.a(new_n20741), .b(new_n20740), .O(new_n20742));
  nor2 g20549(.a(new_n20564), .b(new_n20434), .O(new_n20743));
  inv1 g20550(.a(new_n20743), .O(new_n20744));
  nor2 g20551(.a(new_n20744), .b(new_n20742), .O(new_n20745));
  inv1 g20552(.a(new_n20742), .O(new_n20746));
  nor2 g20553(.a(new_n20743), .b(new_n20746), .O(new_n20747));
  nor2 g20554(.a(new_n20747), .b(new_n20745), .O(new_n20748));
  inv1 g20555(.a(new_n20748), .O(new_n20749));
  nor2 g20556(.a(new_n20574), .b(new_n20568), .O(new_n20750));
  nor2 g20557(.a(new_n20750), .b(new_n20749), .O(new_n20751));
  inv1 g20558(.a(new_n20750), .O(new_n20752));
  nor2 g20559(.a(new_n20752), .b(new_n20748), .O(new_n20753));
  nor2 g20560(.a(new_n20753), .b(new_n20751), .O(\asquared[97] ));
  nor2 g20561(.a(new_n20740), .b(new_n20735), .O(new_n20755));
  nor2 g20562(.a(new_n20729), .b(new_n20723), .O(new_n20756));
  inv1 g20563(.a(new_n20756), .O(new_n20757));
  nor2 g20564(.a(new_n10895), .b(new_n3870), .O(new_n20758));
  inv1 g20565(.a(new_n20758), .O(new_n20759));
  nor2 g20566(.a(new_n20716), .b(new_n20708), .O(new_n20760));
  inv1 g20567(.a(new_n20760), .O(new_n20761));
  nor2 g20568(.a(new_n20761), .b(new_n20759), .O(new_n20762));
  nor2 g20569(.a(new_n20760), .b(new_n20758), .O(new_n20763));
  nor2 g20570(.a(new_n20763), .b(new_n20762), .O(new_n20764));
  nor2 g20571(.a(new_n20697), .b(new_n20689), .O(new_n20765));
  nor2 g20572(.a(new_n20765), .b(new_n20764), .O(new_n20766));
  inv1 g20573(.a(new_n20764), .O(new_n20767));
  inv1 g20574(.a(new_n20765), .O(new_n20768));
  nor2 g20575(.a(new_n20768), .b(new_n20767), .O(new_n20769));
  nor2 g20576(.a(new_n20769), .b(new_n20766), .O(new_n20770));
  inv1 g20577(.a(new_n20770), .O(new_n20771));
  nor2 g20578(.a(new_n20718), .b(new_n20699), .O(new_n20772));
  inv1 g20579(.a(new_n20772), .O(new_n20773));
  nor2 g20580(.a(new_n20659), .b(new_n20653), .O(new_n20774));
  inv1 g20581(.a(new_n20774), .O(new_n20775));
  nor2 g20582(.a(new_n20775), .b(new_n20773), .O(new_n20776));
  nor2 g20583(.a(new_n20774), .b(new_n20772), .O(new_n20777));
  nor2 g20584(.a(new_n20777), .b(new_n20776), .O(new_n20778));
  inv1 g20585(.a(new_n20778), .O(new_n20779));
  nor2 g20586(.a(new_n20779), .b(new_n20771), .O(new_n20780));
  nor2 g20587(.a(new_n20778), .b(new_n20770), .O(new_n20781));
  nor2 g20588(.a(new_n20781), .b(new_n20780), .O(new_n20782));
  inv1 g20589(.a(new_n20782), .O(new_n20783));
  nor2 g20590(.a(new_n20590), .b(new_n20584), .O(new_n20784));
  inv1 g20591(.a(new_n20784), .O(new_n20785));
  nor2 g20592(.a(new_n7537), .b(new_n6274), .O(new_n20786));
  nor2 g20593(.a(new_n20786), .b(new_n20710), .O(new_n20787));
  nor2 g20594(.a(new_n7537), .b(new_n6570), .O(new_n20788));
  inv1 g20595(.a(new_n20788), .O(new_n20789));
  nor2 g20596(.a(new_n20789), .b(new_n20489), .O(new_n20790));
  nor2 g20597(.a(new_n20790), .b(new_n20787), .O(new_n20791));
  nor2 g20598(.a(new_n20791), .b(new_n20538), .O(new_n20792));
  inv1 g20599(.a(new_n20791), .O(new_n20793));
  nor2 g20600(.a(new_n20793), .b(new_n20537), .O(new_n20794));
  nor2 g20601(.a(new_n20794), .b(new_n20792), .O(new_n20795));
  nor2 g20602(.a(new_n6958), .b(\a[48] ), .O(new_n20796));
  nor2 g20603(.a(new_n20796), .b(new_n20617), .O(new_n20797));
  inv1 g20604(.a(new_n20796), .O(new_n20798));
  nor2 g20605(.a(new_n20798), .b(new_n20616), .O(new_n20799));
  nor2 g20606(.a(new_n20799), .b(new_n20797), .O(new_n20800));
  nor2 g20607(.a(new_n20800), .b(new_n20795), .O(new_n20801));
  inv1 g20608(.a(new_n20795), .O(new_n20802));
  inv1 g20609(.a(new_n20800), .O(new_n20803));
  nor2 g20610(.a(new_n20803), .b(new_n20802), .O(new_n20804));
  nor2 g20611(.a(new_n20804), .b(new_n20801), .O(new_n20805));
  nor2 g20612(.a(new_n20805), .b(new_n20785), .O(new_n20806));
  inv1 g20613(.a(new_n20805), .O(new_n20807));
  nor2 g20614(.a(new_n20807), .b(new_n20784), .O(new_n20808));
  nor2 g20615(.a(new_n20808), .b(new_n20806), .O(new_n20809));
  inv1 g20616(.a(new_n20809), .O(new_n20810));
  nor2 g20617(.a(new_n20685), .b(new_n20679), .O(new_n20811));
  nor2 g20618(.a(new_n20621), .b(new_n20614), .O(new_n20812));
  nor2 g20619(.a(new_n20812), .b(new_n20811), .O(new_n20813));
  inv1 g20620(.a(new_n20811), .O(new_n20814));
  inv1 g20621(.a(new_n20812), .O(new_n20815));
  nor2 g20622(.a(new_n20815), .b(new_n20814), .O(new_n20816));
  nor2 g20623(.a(new_n20816), .b(new_n20813), .O(new_n20817));
  nor2 g20624(.a(new_n20636), .b(new_n20629), .O(new_n20818));
  nor2 g20625(.a(new_n20818), .b(new_n20817), .O(new_n20819));
  inv1 g20626(.a(new_n20817), .O(new_n20820));
  inv1 g20627(.a(new_n20818), .O(new_n20821));
  nor2 g20628(.a(new_n20821), .b(new_n20820), .O(new_n20822));
  nor2 g20629(.a(new_n20822), .b(new_n20819), .O(new_n20823));
  nor2 g20630(.a(new_n20645), .b(new_n20638), .O(new_n20824));
  inv1 g20631(.a(new_n20824), .O(new_n20825));
  nor2 g20632(.a(new_n20825), .b(new_n20823), .O(new_n20826));
  inv1 g20633(.a(new_n20823), .O(new_n20827));
  nor2 g20634(.a(new_n20824), .b(new_n20827), .O(new_n20828));
  nor2 g20635(.a(new_n20828), .b(new_n20826), .O(new_n20829));
  inv1 g20636(.a(new_n20829), .O(new_n20830));
  nor2 g20637(.a(new_n20830), .b(new_n20810), .O(new_n20831));
  nor2 g20638(.a(new_n20829), .b(new_n20809), .O(new_n20832));
  nor2 g20639(.a(new_n20832), .b(new_n20831), .O(new_n20833));
  inv1 g20640(.a(new_n20833), .O(new_n20834));
  nor2 g20641(.a(new_n20834), .b(new_n20783), .O(new_n20835));
  nor2 g20642(.a(new_n20833), .b(new_n20782), .O(new_n20836));
  nor2 g20643(.a(new_n20836), .b(new_n20835), .O(new_n20837));
  nor2 g20644(.a(new_n20837), .b(new_n20757), .O(new_n20838));
  inv1 g20645(.a(new_n20837), .O(new_n20839));
  nor2 g20646(.a(new_n20839), .b(new_n20756), .O(new_n20840));
  nor2 g20647(.a(new_n20840), .b(new_n20838), .O(new_n20841));
  inv1 g20648(.a(new_n20841), .O(new_n20842));
  nor2 g20649(.a(new_n20672), .b(new_n20605), .O(new_n20843));
  inv1 g20650(.a(new_n20843), .O(new_n20844));
  nor2 g20651(.a(new_n20668), .b(new_n20665), .O(new_n20845));
  nor2 g20652(.a(new_n20601), .b(new_n20598), .O(new_n20846));
  nor2 g20653(.a(new_n8026), .b(new_n5971), .O(new_n20847));
  nor2 g20654(.a(new_n8170), .b(new_n5796), .O(new_n20848));
  nor2 g20655(.a(new_n20848), .b(new_n20847), .O(new_n20849));
  nor2 g20656(.a(new_n8170), .b(new_n5971), .O(new_n20850));
  inv1 g20657(.a(new_n20850), .O(new_n20851));
  nor2 g20658(.a(new_n20851), .b(new_n20475), .O(new_n20852));
  nor2 g20659(.a(new_n20852), .b(new_n20849), .O(new_n20853));
  nor2 g20660(.a(new_n20853), .b(new_n20631), .O(new_n20854));
  inv1 g20661(.a(new_n20853), .O(new_n20855));
  nor2 g20662(.a(new_n20855), .b(new_n20630), .O(new_n20856));
  nor2 g20663(.a(new_n20856), .b(new_n20854), .O(new_n20857));
  nor2 g20664(.a(new_n10468), .b(new_n4093), .O(new_n20858));
  inv1 g20665(.a(new_n20858), .O(new_n20859));
  nor2 g20666(.a(new_n10320), .b(new_n4366), .O(new_n20860));
  nor2 g20667(.a(new_n20860), .b(new_n20691), .O(new_n20861));
  inv1 g20668(.a(new_n20688), .O(new_n20862));
  nor2 g20669(.a(new_n10320), .b(new_n4425), .O(new_n20863));
  inv1 g20670(.a(new_n20863), .O(new_n20864));
  nor2 g20671(.a(new_n20864), .b(new_n20862), .O(new_n20865));
  nor2 g20672(.a(new_n20865), .b(new_n20861), .O(new_n20866));
  nor2 g20673(.a(new_n20866), .b(new_n20859), .O(new_n20867));
  inv1 g20674(.a(new_n20866), .O(new_n20868));
  nor2 g20675(.a(new_n20868), .b(new_n20858), .O(new_n20869));
  nor2 g20676(.a(new_n20869), .b(new_n20867), .O(new_n20870));
  nor2 g20677(.a(new_n9156), .b(new_n4954), .O(new_n20871));
  inv1 g20678(.a(new_n20871), .O(new_n20872));
  nor2 g20679(.a(new_n8946), .b(new_n5178), .O(new_n20873));
  nor2 g20680(.a(new_n20873), .b(new_n20522), .O(new_n20874));
  inv1 g20681(.a(new_n20873), .O(new_n20875));
  nor2 g20682(.a(new_n20875), .b(new_n20523), .O(new_n20876));
  nor2 g20683(.a(new_n20876), .b(new_n20874), .O(new_n20877));
  nor2 g20684(.a(new_n20877), .b(new_n20872), .O(new_n20878));
  inv1 g20685(.a(new_n20877), .O(new_n20879));
  nor2 g20686(.a(new_n20879), .b(new_n20871), .O(new_n20880));
  nor2 g20687(.a(new_n20880), .b(new_n20878), .O(new_n20881));
  nor2 g20688(.a(new_n20881), .b(new_n20870), .O(new_n20882));
  inv1 g20689(.a(new_n20870), .O(new_n20883));
  inv1 g20690(.a(new_n20881), .O(new_n20884));
  nor2 g20691(.a(new_n20884), .b(new_n20883), .O(new_n20885));
  nor2 g20692(.a(new_n20885), .b(new_n20882), .O(new_n20886));
  inv1 g20693(.a(new_n20886), .O(new_n20887));
  nor2 g20694(.a(new_n20887), .b(new_n20857), .O(new_n20888));
  inv1 g20695(.a(new_n20857), .O(new_n20889));
  nor2 g20696(.a(new_n20886), .b(new_n20889), .O(new_n20890));
  nor2 g20697(.a(new_n20890), .b(new_n20888), .O(new_n20891));
  inv1 g20698(.a(new_n20891), .O(new_n20892));
  nor2 g20699(.a(new_n20892), .b(new_n20846), .O(new_n20893));
  inv1 g20700(.a(new_n20846), .O(new_n20894));
  nor2 g20701(.a(new_n20891), .b(new_n20894), .O(new_n20895));
  nor2 g20702(.a(new_n20895), .b(new_n20893), .O(new_n20896));
  inv1 g20703(.a(new_n20896), .O(new_n20897));
  nor2 g20704(.a(new_n20897), .b(new_n20845), .O(new_n20898));
  inv1 g20705(.a(new_n20845), .O(new_n20899));
  nor2 g20706(.a(new_n20896), .b(new_n20899), .O(new_n20900));
  nor2 g20707(.a(new_n20900), .b(new_n20898), .O(new_n20901));
  nor2 g20708(.a(new_n20901), .b(new_n20844), .O(new_n20902));
  inv1 g20709(.a(new_n20901), .O(new_n20903));
  nor2 g20710(.a(new_n20903), .b(new_n20843), .O(new_n20904));
  nor2 g20711(.a(new_n20904), .b(new_n20902), .O(new_n20905));
  inv1 g20712(.a(new_n20905), .O(new_n20906));
  nor2 g20713(.a(new_n20906), .b(new_n20842), .O(new_n20907));
  nor2 g20714(.a(new_n20905), .b(new_n20841), .O(new_n20908));
  nor2 g20715(.a(new_n20908), .b(new_n20907), .O(new_n20909));
  inv1 g20716(.a(new_n20909), .O(new_n20910));
  nor2 g20717(.a(new_n20910), .b(new_n20755), .O(new_n20911));
  inv1 g20718(.a(new_n20755), .O(new_n20912));
  nor2 g20719(.a(new_n20909), .b(new_n20912), .O(new_n20913));
  nor2 g20720(.a(new_n20913), .b(new_n20911), .O(new_n20914));
  inv1 g20721(.a(new_n20914), .O(new_n20915));
  nor2 g20722(.a(new_n20751), .b(new_n20747), .O(new_n20916));
  inv1 g20723(.a(new_n20916), .O(new_n20917));
  nor2 g20724(.a(new_n20917), .b(new_n20915), .O(new_n20918));
  nor2 g20725(.a(new_n20916), .b(new_n20914), .O(new_n20919));
  nor2 g20726(.a(new_n20919), .b(new_n20918), .O(new_n20920));
  inv1 g20727(.a(new_n20920), .O(\asquared[98] ));
  nor2 g20728(.a(new_n20907), .b(new_n20904), .O(new_n20922));
  inv1 g20729(.a(new_n20922), .O(new_n20923));
  nor2 g20730(.a(new_n20898), .b(new_n20893), .O(new_n20924));
  nor2 g20731(.a(new_n20822), .b(new_n20816), .O(new_n20925));
  inv1 g20732(.a(new_n20925), .O(new_n20926));
  nor2 g20733(.a(new_n20769), .b(new_n20762), .O(new_n20927));
  inv1 g20734(.a(new_n20927), .O(new_n20928));
  nor2 g20735(.a(new_n20928), .b(new_n20926), .O(new_n20929));
  nor2 g20736(.a(new_n20927), .b(new_n20925), .O(new_n20930));
  nor2 g20737(.a(new_n20930), .b(new_n20929), .O(new_n20931));
  nor2 g20738(.a(new_n20888), .b(new_n20882), .O(new_n20932));
  inv1 g20739(.a(new_n20932), .O(new_n20933));
  nor2 g20740(.a(new_n20933), .b(new_n20931), .O(new_n20934));
  inv1 g20741(.a(new_n20931), .O(new_n20935));
  nor2 g20742(.a(new_n20932), .b(new_n20935), .O(new_n20936));
  nor2 g20743(.a(new_n20936), .b(new_n20934), .O(new_n20937));
  inv1 g20744(.a(new_n20937), .O(new_n20938));
  nor2 g20745(.a(new_n20880), .b(new_n20874), .O(new_n20939));
  nor2 g20746(.a(new_n20869), .b(new_n20861), .O(new_n20940));
  nor2 g20747(.a(new_n20940), .b(new_n20939), .O(new_n20941));
  inv1 g20748(.a(new_n20939), .O(new_n20942));
  inv1 g20749(.a(new_n20940), .O(new_n20943));
  nor2 g20750(.a(new_n20943), .b(new_n20942), .O(new_n20944));
  nor2 g20751(.a(new_n20944), .b(new_n20941), .O(new_n20945));
  nor2 g20752(.a(new_n20856), .b(new_n20849), .O(new_n20946));
  nor2 g20753(.a(new_n20946), .b(new_n20945), .O(new_n20947));
  inv1 g20754(.a(new_n20945), .O(new_n20948));
  inv1 g20755(.a(new_n20946), .O(new_n20949));
  nor2 g20756(.a(new_n20949), .b(new_n20948), .O(new_n20950));
  nor2 g20757(.a(new_n20950), .b(new_n20947), .O(new_n20951));
  nor2 g20758(.a(new_n20808), .b(new_n20801), .O(new_n20952));
  inv1 g20759(.a(new_n20952), .O(new_n20953));
  nor2 g20760(.a(new_n20953), .b(new_n20951), .O(new_n20954));
  inv1 g20761(.a(new_n20951), .O(new_n20955));
  nor2 g20762(.a(new_n20952), .b(new_n20955), .O(new_n20956));
  nor2 g20763(.a(new_n20956), .b(new_n20954), .O(new_n20957));
  inv1 g20764(.a(new_n20957), .O(new_n20958));
  nor2 g20765(.a(new_n10895), .b(new_n4093), .O(new_n20959));
  nor2 g20766(.a(new_n20959), .b(new_n14406), .O(new_n20960));
  nor2 g20767(.a(new_n11186), .b(new_n4093), .O(new_n20961));
  inv1 g20768(.a(new_n20961), .O(new_n20962));
  nor2 g20769(.a(new_n20962), .b(new_n20759), .O(new_n20963));
  nor2 g20770(.a(new_n20963), .b(new_n20960), .O(new_n20964));
  inv1 g20771(.a(new_n20964), .O(new_n20965));
  nor2 g20772(.a(new_n20799), .b(new_n6958), .O(new_n20966));
  inv1 g20773(.a(new_n20966), .O(new_n20967));
  nor2 g20774(.a(new_n20967), .b(new_n20965), .O(new_n20968));
  nor2 g20775(.a(new_n20966), .b(new_n20964), .O(new_n20969));
  nor2 g20776(.a(new_n20969), .b(new_n20968), .O(new_n20970));
  inv1 g20777(.a(new_n20970), .O(new_n20971));
  nor2 g20778(.a(new_n9873), .b(new_n4682), .O(new_n20972));
  nor2 g20779(.a(new_n20972), .b(new_n20863), .O(new_n20973));
  nor2 g20780(.a(new_n20692), .b(new_n20681), .O(new_n20974));
  nor2 g20781(.a(new_n20974), .b(new_n20973), .O(new_n20975));
  inv1 g20782(.a(new_n20975), .O(new_n20976));
  nor2 g20783(.a(new_n20976), .b(new_n20850), .O(new_n20977));
  nor2 g20784(.a(new_n20975), .b(new_n20851), .O(new_n20978));
  nor2 g20785(.a(new_n20978), .b(new_n20977), .O(new_n20979));
  nor2 g20786(.a(new_n8026), .b(new_n6274), .O(new_n20980));
  inv1 g20787(.a(new_n20980), .O(new_n20981));
  nor2 g20788(.a(new_n7294), .b(new_n6893), .O(new_n20982));
  nor2 g20789(.a(new_n20982), .b(new_n20788), .O(new_n20983));
  nor2 g20790(.a(new_n7537), .b(new_n6893), .O(new_n20984));
  inv1 g20791(.a(new_n20984), .O(new_n20985));
  nor2 g20792(.a(new_n20985), .b(new_n20711), .O(new_n20986));
  nor2 g20793(.a(new_n20986), .b(new_n20983), .O(new_n20987));
  nor2 g20794(.a(new_n20987), .b(new_n20981), .O(new_n20988));
  inv1 g20795(.a(new_n20987), .O(new_n20989));
  nor2 g20796(.a(new_n20989), .b(new_n20980), .O(new_n20990));
  nor2 g20797(.a(new_n20990), .b(new_n20988), .O(new_n20991));
  nor2 g20798(.a(new_n20991), .b(new_n20979), .O(new_n20992));
  inv1 g20799(.a(new_n20979), .O(new_n20993));
  inv1 g20800(.a(new_n20991), .O(new_n20994));
  nor2 g20801(.a(new_n20994), .b(new_n20993), .O(new_n20995));
  nor2 g20802(.a(new_n20995), .b(new_n20992), .O(new_n20996));
  inv1 g20803(.a(new_n20996), .O(new_n20997));
  nor2 g20804(.a(new_n20997), .b(new_n20971), .O(new_n20998));
  nor2 g20805(.a(new_n20996), .b(new_n20970), .O(new_n20999));
  nor2 g20806(.a(new_n20999), .b(new_n20998), .O(new_n21000));
  inv1 g20807(.a(new_n21000), .O(new_n21001));
  nor2 g20808(.a(new_n21001), .b(new_n20958), .O(new_n21002));
  nor2 g20809(.a(new_n21000), .b(new_n20957), .O(new_n21003));
  nor2 g20810(.a(new_n21003), .b(new_n21002), .O(new_n21004));
  inv1 g20811(.a(new_n21004), .O(new_n21005));
  nor2 g20812(.a(new_n21005), .b(new_n20938), .O(new_n21006));
  nor2 g20813(.a(new_n21004), .b(new_n20937), .O(new_n21007));
  nor2 g20814(.a(new_n21007), .b(new_n21006), .O(new_n21008));
  inv1 g20815(.a(new_n21008), .O(new_n21009));
  nor2 g20816(.a(new_n21009), .b(new_n20924), .O(new_n21010));
  inv1 g20817(.a(new_n20924), .O(new_n21011));
  nor2 g20818(.a(new_n21008), .b(new_n21011), .O(new_n21012));
  nor2 g20819(.a(new_n21012), .b(new_n21010), .O(new_n21013));
  inv1 g20820(.a(new_n21013), .O(new_n21014));
  nor2 g20821(.a(new_n20840), .b(new_n20835), .O(new_n21015));
  nor2 g20822(.a(new_n20831), .b(new_n20828), .O(new_n21016));
  nor2 g20823(.a(new_n20780), .b(new_n20777), .O(new_n21017));
  nor2 g20824(.a(new_n8946), .b(new_n5393), .O(new_n21018));
  nor2 g20825(.a(new_n8476), .b(new_n5796), .O(new_n21019));
  nor2 g20826(.a(new_n21019), .b(new_n21018), .O(new_n21020));
  nor2 g20827(.a(new_n8946), .b(new_n5796), .O(new_n21021));
  inv1 g20828(.a(new_n21021), .O(new_n21022));
  nor2 g20829(.a(new_n21022), .b(new_n20631), .O(new_n21023));
  nor2 g20830(.a(new_n21023), .b(new_n21020), .O(new_n21024));
  nor2 g20831(.a(new_n11596), .b(new_n3722), .O(new_n21025));
  nor2 g20832(.a(new_n21025), .b(new_n21024), .O(new_n21026));
  inv1 g20833(.a(new_n21024), .O(new_n21027));
  inv1 g20834(.a(new_n21025), .O(new_n21028));
  nor2 g20835(.a(new_n21028), .b(new_n21027), .O(new_n21029));
  nor2 g20836(.a(new_n21029), .b(new_n21026), .O(new_n21030));
  inv1 g20837(.a(new_n21030), .O(new_n21031));
  nor2 g20838(.a(new_n20794), .b(new_n20787), .O(new_n21032));
  inv1 g20839(.a(new_n21032), .O(new_n21033));
  nor2 g20840(.a(new_n21033), .b(new_n21031), .O(new_n21034));
  nor2 g20841(.a(new_n21032), .b(new_n21030), .O(new_n21035));
  nor2 g20842(.a(new_n21035), .b(new_n21034), .O(new_n21036));
  inv1 g20843(.a(new_n21036), .O(new_n21037));
  nor2 g20844(.a(new_n10468), .b(new_n4366), .O(new_n21038));
  inv1 g20845(.a(new_n21038), .O(new_n21039));
  nor2 g20846(.a(new_n9156), .b(new_n5178), .O(new_n21040));
  nor2 g20847(.a(new_n9658), .b(new_n4954), .O(new_n21041));
  nor2 g20848(.a(new_n21041), .b(new_n21040), .O(new_n21042));
  nor2 g20849(.a(new_n9658), .b(new_n5178), .O(new_n21043));
  inv1 g20850(.a(new_n21043), .O(new_n21044));
  nor2 g20851(.a(new_n21044), .b(new_n20872), .O(new_n21045));
  nor2 g20852(.a(new_n21045), .b(new_n21042), .O(new_n21046));
  nor2 g20853(.a(new_n21046), .b(new_n21039), .O(new_n21047));
  inv1 g20854(.a(new_n21046), .O(new_n21048));
  nor2 g20855(.a(new_n21048), .b(new_n21038), .O(new_n21049));
  nor2 g20856(.a(new_n21049), .b(new_n21047), .O(new_n21050));
  nor2 g20857(.a(new_n21050), .b(new_n21037), .O(new_n21051));
  inv1 g20858(.a(new_n21050), .O(new_n21052));
  nor2 g20859(.a(new_n21052), .b(new_n21036), .O(new_n21053));
  nor2 g20860(.a(new_n21053), .b(new_n21051), .O(new_n21054));
  inv1 g20861(.a(new_n21054), .O(new_n21055));
  nor2 g20862(.a(new_n21055), .b(new_n21017), .O(new_n21056));
  inv1 g20863(.a(new_n21017), .O(new_n21057));
  nor2 g20864(.a(new_n21054), .b(new_n21057), .O(new_n21058));
  nor2 g20865(.a(new_n21058), .b(new_n21056), .O(new_n21059));
  inv1 g20866(.a(new_n21059), .O(new_n21060));
  nor2 g20867(.a(new_n21060), .b(new_n21016), .O(new_n21061));
  inv1 g20868(.a(new_n21016), .O(new_n21062));
  nor2 g20869(.a(new_n21059), .b(new_n21062), .O(new_n21063));
  nor2 g20870(.a(new_n21063), .b(new_n21061), .O(new_n21064));
  inv1 g20871(.a(new_n21064), .O(new_n21065));
  nor2 g20872(.a(new_n21065), .b(new_n21015), .O(new_n21066));
  inv1 g20873(.a(new_n21015), .O(new_n21067));
  nor2 g20874(.a(new_n21064), .b(new_n21067), .O(new_n21068));
  nor2 g20875(.a(new_n21068), .b(new_n21066), .O(new_n21069));
  inv1 g20876(.a(new_n21069), .O(new_n21070));
  nor2 g20877(.a(new_n21070), .b(new_n21014), .O(new_n21071));
  nor2 g20878(.a(new_n21069), .b(new_n21013), .O(new_n21072));
  nor2 g20879(.a(new_n21072), .b(new_n21071), .O(new_n21073));
  nor2 g20880(.a(new_n21073), .b(new_n20923), .O(new_n21074));
  inv1 g20881(.a(new_n21073), .O(new_n21075));
  nor2 g20882(.a(new_n21075), .b(new_n20922), .O(new_n21076));
  nor2 g20883(.a(new_n21076), .b(new_n21074), .O(new_n21077));
  inv1 g20884(.a(new_n21077), .O(new_n21078));
  nor2 g20885(.a(new_n20916), .b(new_n20913), .O(new_n21079));
  nor2 g20886(.a(new_n21079), .b(new_n20911), .O(new_n21080));
  nor2 g20887(.a(new_n21080), .b(new_n21078), .O(new_n21081));
  inv1 g20888(.a(new_n21080), .O(new_n21082));
  nor2 g20889(.a(new_n21082), .b(new_n21077), .O(new_n21083));
  nor2 g20890(.a(new_n21083), .b(new_n21081), .O(\asquared[99] ));
  nor2 g20891(.a(new_n21071), .b(new_n21066), .O(new_n21085));
  nor2 g20892(.a(new_n21061), .b(new_n21056), .O(new_n21086));
  nor2 g20893(.a(new_n21051), .b(new_n21034), .O(new_n21087));
  inv1 g20894(.a(new_n21087), .O(new_n21088));
  nor2 g20895(.a(new_n20950), .b(new_n20944), .O(new_n21089));
  nor2 g20896(.a(new_n7294), .b(\a[49] ), .O(new_n21090));
  nor2 g20897(.a(new_n21090), .b(new_n20962), .O(new_n21091));
  inv1 g20898(.a(new_n21090), .O(new_n21092));
  nor2 g20899(.a(new_n21092), .b(new_n20961), .O(new_n21093));
  nor2 g20900(.a(new_n21093), .b(new_n21091), .O(new_n21094));
  nor2 g20901(.a(new_n21094), .b(new_n21089), .O(new_n21095));
  inv1 g20902(.a(new_n21089), .O(new_n21096));
  inv1 g20903(.a(new_n21094), .O(new_n21097));
  nor2 g20904(.a(new_n21097), .b(new_n21096), .O(new_n21098));
  nor2 g20905(.a(new_n21098), .b(new_n21095), .O(new_n21099));
  nor2 g20906(.a(new_n21099), .b(new_n21088), .O(new_n21100));
  inv1 g20907(.a(new_n21099), .O(new_n21101));
  nor2 g20908(.a(new_n21101), .b(new_n21087), .O(new_n21102));
  nor2 g20909(.a(new_n21102), .b(new_n21100), .O(new_n21103));
  inv1 g20910(.a(new_n21103), .O(new_n21104));
  nor2 g20911(.a(new_n20990), .b(new_n20983), .O(new_n21105));
  nor2 g20912(.a(new_n20977), .b(new_n20973), .O(new_n21106));
  nor2 g20913(.a(new_n21106), .b(new_n21105), .O(new_n21107));
  inv1 g20914(.a(new_n21105), .O(new_n21108));
  inv1 g20915(.a(new_n21106), .O(new_n21109));
  nor2 g20916(.a(new_n21109), .b(new_n21108), .O(new_n21110));
  nor2 g20917(.a(new_n21110), .b(new_n21107), .O(new_n21111));
  nor2 g20918(.a(new_n21029), .b(new_n21023), .O(new_n21112));
  inv1 g20919(.a(new_n21112), .O(new_n21113));
  nor2 g20920(.a(new_n21113), .b(new_n21111), .O(new_n21114));
  inv1 g20921(.a(new_n21111), .O(new_n21115));
  nor2 g20922(.a(new_n21112), .b(new_n21115), .O(new_n21116));
  nor2 g20923(.a(new_n21116), .b(new_n21114), .O(new_n21117));
  inv1 g20924(.a(new_n21117), .O(new_n21118));
  nor2 g20925(.a(new_n20998), .b(new_n20992), .O(new_n21119));
  nor2 g20926(.a(new_n21119), .b(new_n21118), .O(new_n21120));
  inv1 g20927(.a(new_n21119), .O(new_n21121));
  nor2 g20928(.a(new_n21121), .b(new_n21117), .O(new_n21122));
  nor2 g20929(.a(new_n21122), .b(new_n21120), .O(new_n21123));
  inv1 g20930(.a(new_n21123), .O(new_n21124));
  nor2 g20931(.a(new_n20968), .b(new_n20963), .O(new_n21125));
  inv1 g20932(.a(new_n21125), .O(new_n21126));
  nor2 g20933(.a(new_n21049), .b(new_n21042), .O(new_n21127));
  nor2 g20934(.a(new_n21127), .b(new_n21126), .O(new_n21128));
  inv1 g20935(.a(new_n21127), .O(new_n21129));
  nor2 g20936(.a(new_n21129), .b(new_n21125), .O(new_n21130));
  nor2 g20937(.a(new_n21130), .b(new_n21128), .O(new_n21131));
  inv1 g20938(.a(new_n21131), .O(new_n21132));
  nor2 g20939(.a(new_n11596), .b(new_n3870), .O(new_n21133));
  inv1 g20940(.a(new_n21133), .O(new_n21134));
  nor2 g20941(.a(new_n10468), .b(new_n4425), .O(new_n21135));
  nor2 g20942(.a(new_n10895), .b(new_n4366), .O(new_n21136));
  nor2 g20943(.a(new_n21136), .b(new_n21135), .O(new_n21137));
  nor2 g20944(.a(new_n10895), .b(new_n4425), .O(new_n21138));
  inv1 g20945(.a(new_n21138), .O(new_n21139));
  nor2 g20946(.a(new_n21139), .b(new_n21039), .O(new_n21140));
  nor2 g20947(.a(new_n21140), .b(new_n21137), .O(new_n21141));
  nor2 g20948(.a(new_n21141), .b(new_n21134), .O(new_n21142));
  inv1 g20949(.a(new_n21141), .O(new_n21143));
  nor2 g20950(.a(new_n21143), .b(new_n21133), .O(new_n21144));
  nor2 g20951(.a(new_n21144), .b(new_n21142), .O(new_n21145));
  nor2 g20952(.a(new_n21145), .b(new_n21132), .O(new_n21146));
  inv1 g20953(.a(new_n21145), .O(new_n21147));
  nor2 g20954(.a(new_n21147), .b(new_n21131), .O(new_n21148));
  nor2 g20955(.a(new_n21148), .b(new_n21146), .O(new_n21149));
  inv1 g20956(.a(new_n21149), .O(new_n21150));
  nor2 g20957(.a(new_n21150), .b(new_n21124), .O(new_n21151));
  nor2 g20958(.a(new_n21149), .b(new_n21123), .O(new_n21152));
  nor2 g20959(.a(new_n21152), .b(new_n21151), .O(new_n21153));
  inv1 g20960(.a(new_n21153), .O(new_n21154));
  nor2 g20961(.a(new_n21154), .b(new_n21104), .O(new_n21155));
  nor2 g20962(.a(new_n21153), .b(new_n21103), .O(new_n21156));
  nor2 g20963(.a(new_n21156), .b(new_n21155), .O(new_n21157));
  inv1 g20964(.a(new_n21157), .O(new_n21158));
  nor2 g20965(.a(new_n21158), .b(new_n21086), .O(new_n21159));
  inv1 g20966(.a(new_n21086), .O(new_n21160));
  nor2 g20967(.a(new_n21157), .b(new_n21160), .O(new_n21161));
  nor2 g20968(.a(new_n21161), .b(new_n21159), .O(new_n21162));
  inv1 g20969(.a(new_n21162), .O(new_n21163));
  nor2 g20970(.a(new_n20936), .b(new_n20930), .O(new_n21164));
  inv1 g20971(.a(new_n21164), .O(new_n21165));
  nor2 g20972(.a(new_n9156), .b(new_n5393), .O(new_n21166));
  nor2 g20973(.a(new_n21166), .b(new_n21043), .O(new_n21167));
  inv1 g20974(.a(new_n21040), .O(new_n21168));
  nor2 g20975(.a(new_n9658), .b(new_n5393), .O(new_n21169));
  inv1 g20976(.a(new_n21169), .O(new_n21170));
  nor2 g20977(.a(new_n21170), .b(new_n21168), .O(new_n21171));
  nor2 g20978(.a(new_n21171), .b(new_n21167), .O(new_n21172));
  nor2 g20979(.a(new_n21172), .b(new_n20985), .O(new_n21173));
  inv1 g20980(.a(new_n21172), .O(new_n21174));
  nor2 g20981(.a(new_n21174), .b(new_n20984), .O(new_n21175));
  nor2 g20982(.a(new_n21175), .b(new_n21173), .O(new_n21176));
  inv1 g20983(.a(new_n21176), .O(new_n21177));
  nor2 g20984(.a(new_n8476), .b(new_n5971), .O(new_n21178));
  inv1 g20985(.a(new_n21178), .O(new_n21179));
  nor2 g20986(.a(new_n8026), .b(new_n6570), .O(new_n21180));
  nor2 g20987(.a(new_n8170), .b(new_n6274), .O(new_n21181));
  nor2 g20988(.a(new_n21181), .b(new_n21180), .O(new_n21182));
  nor2 g20989(.a(new_n8170), .b(new_n6570), .O(new_n21183));
  inv1 g20990(.a(new_n21183), .O(new_n21184));
  nor2 g20991(.a(new_n21184), .b(new_n20981), .O(new_n21185));
  nor2 g20992(.a(new_n21185), .b(new_n21182), .O(new_n21186));
  nor2 g20993(.a(new_n21186), .b(new_n21179), .O(new_n21187));
  inv1 g20994(.a(new_n21186), .O(new_n21188));
  nor2 g20995(.a(new_n21188), .b(new_n21178), .O(new_n21189));
  nor2 g20996(.a(new_n21189), .b(new_n21187), .O(new_n21190));
  nor2 g20997(.a(new_n9873), .b(new_n4954), .O(new_n21191));
  nor2 g20998(.a(new_n21191), .b(new_n21021), .O(new_n21192));
  inv1 g20999(.a(new_n21191), .O(new_n21193));
  nor2 g21000(.a(new_n21193), .b(new_n21022), .O(new_n21194));
  nor2 g21001(.a(new_n21194), .b(new_n21192), .O(new_n21195));
  nor2 g21002(.a(new_n21195), .b(new_n20681), .O(new_n21196));
  inv1 g21003(.a(new_n21195), .O(new_n21197));
  nor2 g21004(.a(new_n21197), .b(new_n20680), .O(new_n21198));
  nor2 g21005(.a(new_n21198), .b(new_n21196), .O(new_n21199));
  nor2 g21006(.a(new_n21199), .b(new_n21190), .O(new_n21200));
  inv1 g21007(.a(new_n21190), .O(new_n21201));
  inv1 g21008(.a(new_n21199), .O(new_n21202));
  nor2 g21009(.a(new_n21202), .b(new_n21201), .O(new_n21203));
  nor2 g21010(.a(new_n21203), .b(new_n21200), .O(new_n21204));
  nor2 g21011(.a(new_n21204), .b(new_n21177), .O(new_n21205));
  inv1 g21012(.a(new_n21204), .O(new_n21206));
  nor2 g21013(.a(new_n21206), .b(new_n21176), .O(new_n21207));
  nor2 g21014(.a(new_n21207), .b(new_n21205), .O(new_n21208));
  nor2 g21015(.a(new_n21208), .b(new_n21165), .O(new_n21209));
  inv1 g21016(.a(new_n21208), .O(new_n21210));
  nor2 g21017(.a(new_n21210), .b(new_n21164), .O(new_n21211));
  nor2 g21018(.a(new_n21211), .b(new_n21209), .O(new_n21212));
  nor2 g21019(.a(new_n21002), .b(new_n20956), .O(new_n21213));
  inv1 g21020(.a(new_n21213), .O(new_n21214));
  nor2 g21021(.a(new_n21214), .b(new_n21212), .O(new_n21215));
  inv1 g21022(.a(new_n21212), .O(new_n21216));
  nor2 g21023(.a(new_n21213), .b(new_n21216), .O(new_n21217));
  nor2 g21024(.a(new_n21217), .b(new_n21215), .O(new_n21218));
  inv1 g21025(.a(new_n21218), .O(new_n21219));
  nor2 g21026(.a(new_n21010), .b(new_n21006), .O(new_n21220));
  nor2 g21027(.a(new_n21220), .b(new_n21219), .O(new_n21221));
  inv1 g21028(.a(new_n21220), .O(new_n21222));
  nor2 g21029(.a(new_n21222), .b(new_n21218), .O(new_n21223));
  nor2 g21030(.a(new_n21223), .b(new_n21221), .O(new_n21224));
  inv1 g21031(.a(new_n21224), .O(new_n21225));
  nor2 g21032(.a(new_n21225), .b(new_n21163), .O(new_n21226));
  nor2 g21033(.a(new_n21224), .b(new_n21162), .O(new_n21227));
  nor2 g21034(.a(new_n21227), .b(new_n21226), .O(new_n21228));
  inv1 g21035(.a(new_n21228), .O(new_n21229));
  nor2 g21036(.a(new_n21229), .b(new_n21085), .O(new_n21230));
  inv1 g21037(.a(new_n21085), .O(new_n21231));
  nor2 g21038(.a(new_n21228), .b(new_n21231), .O(new_n21232));
  nor2 g21039(.a(new_n21232), .b(new_n21230), .O(new_n21233));
  inv1 g21040(.a(new_n21233), .O(new_n21234));
  nor2 g21041(.a(new_n21081), .b(new_n21076), .O(new_n21235));
  nor2 g21042(.a(new_n21235), .b(new_n21234), .O(new_n21236));
  inv1 g21043(.a(new_n21235), .O(new_n21237));
  nor2 g21044(.a(new_n21237), .b(new_n21233), .O(new_n21238));
  nor2 g21045(.a(new_n21238), .b(new_n21236), .O(\asquared[100] ));
  nor2 g21046(.a(new_n21226), .b(new_n21221), .O(new_n21240));
  nor2 g21047(.a(new_n21116), .b(new_n21110), .O(new_n21241));
  nor2 g21048(.a(new_n7537), .b(new_n6958), .O(new_n21242));
  nor2 g21049(.a(new_n8026), .b(new_n6893), .O(new_n21243));
  nor2 g21050(.a(new_n21243), .b(new_n21242), .O(new_n21244));
  nor2 g21051(.a(new_n8026), .b(new_n6958), .O(new_n21245));
  inv1 g21052(.a(new_n21245), .O(new_n21246));
  nor2 g21053(.a(new_n21246), .b(new_n20985), .O(new_n21247));
  nor2 g21054(.a(new_n21247), .b(new_n21244), .O(new_n21248));
  nor2 g21055(.a(new_n21248), .b(new_n21184), .O(new_n21249));
  inv1 g21056(.a(new_n21248), .O(new_n21250));
  nor2 g21057(.a(new_n21250), .b(new_n21183), .O(new_n21251));
  nor2 g21058(.a(new_n21251), .b(new_n21249), .O(new_n21252));
  nor2 g21059(.a(new_n21252), .b(new_n21241), .O(new_n21253));
  inv1 g21060(.a(new_n21241), .O(new_n21254));
  inv1 g21061(.a(new_n21252), .O(new_n21255));
  nor2 g21062(.a(new_n21255), .b(new_n21254), .O(new_n21256));
  nor2 g21063(.a(new_n21256), .b(new_n21253), .O(new_n21257));
  nor2 g21064(.a(new_n21146), .b(new_n21130), .O(new_n21258));
  inv1 g21065(.a(new_n21258), .O(new_n21259));
  nor2 g21066(.a(new_n21259), .b(new_n21257), .O(new_n21260));
  inv1 g21067(.a(new_n21257), .O(new_n21261));
  nor2 g21068(.a(new_n21258), .b(new_n21261), .O(new_n21262));
  nor2 g21069(.a(new_n21262), .b(new_n21260), .O(new_n21263));
  nor2 g21070(.a(new_n21217), .b(new_n21211), .O(new_n21264));
  inv1 g21071(.a(new_n21264), .O(new_n21265));
  nor2 g21072(.a(new_n21265), .b(new_n21263), .O(new_n21266));
  inv1 g21073(.a(new_n21263), .O(new_n21267));
  nor2 g21074(.a(new_n21264), .b(new_n21267), .O(new_n21268));
  nor2 g21075(.a(new_n21268), .b(new_n21266), .O(new_n21269));
  inv1 g21076(.a(new_n21269), .O(new_n21270));
  nor2 g21077(.a(new_n21144), .b(new_n21137), .O(new_n21271));
  nor2 g21078(.a(new_n21189), .b(new_n21182), .O(new_n21272));
  nor2 g21079(.a(new_n21272), .b(new_n21271), .O(new_n21273));
  inv1 g21080(.a(new_n21271), .O(new_n21274));
  inv1 g21081(.a(new_n21272), .O(new_n21275));
  nor2 g21082(.a(new_n21275), .b(new_n21274), .O(new_n21276));
  nor2 g21083(.a(new_n21276), .b(new_n21273), .O(new_n21277));
  nor2 g21084(.a(new_n21198), .b(new_n21192), .O(new_n21278));
  nor2 g21085(.a(new_n21278), .b(new_n21277), .O(new_n21279));
  inv1 g21086(.a(new_n21277), .O(new_n21280));
  inv1 g21087(.a(new_n21278), .O(new_n21281));
  nor2 g21088(.a(new_n21281), .b(new_n21280), .O(new_n21282));
  nor2 g21089(.a(new_n21282), .b(new_n21279), .O(new_n21283));
  nor2 g21090(.a(new_n21207), .b(new_n21200), .O(new_n21284));
  inv1 g21091(.a(new_n21284), .O(new_n21285));
  nor2 g21092(.a(new_n21285), .b(new_n21283), .O(new_n21286));
  inv1 g21093(.a(new_n21283), .O(new_n21287));
  nor2 g21094(.a(new_n21284), .b(new_n21287), .O(new_n21288));
  nor2 g21095(.a(new_n21288), .b(new_n21286), .O(new_n21289));
  inv1 g21096(.a(new_n21289), .O(new_n21290));
  nor2 g21097(.a(new_n11596), .b(new_n4093), .O(new_n21291));
  inv1 g21098(.a(new_n21291), .O(new_n21292));
  nor2 g21099(.a(new_n21093), .b(new_n7294), .O(new_n21293));
  inv1 g21100(.a(new_n21293), .O(new_n21294));
  nor2 g21101(.a(new_n21294), .b(new_n21292), .O(new_n21295));
  nor2 g21102(.a(new_n21293), .b(new_n21291), .O(new_n21296));
  nor2 g21103(.a(new_n21296), .b(new_n21295), .O(new_n21297));
  nor2 g21104(.a(new_n21175), .b(new_n21167), .O(new_n21298));
  nor2 g21105(.a(new_n21298), .b(new_n21297), .O(new_n21299));
  inv1 g21106(.a(new_n21297), .O(new_n21300));
  inv1 g21107(.a(new_n21298), .O(new_n21301));
  nor2 g21108(.a(new_n21301), .b(new_n21300), .O(new_n21302));
  nor2 g21109(.a(new_n21302), .b(new_n21299), .O(new_n21303));
  inv1 g21110(.a(new_n21303), .O(new_n21304));
  nor2 g21111(.a(new_n21304), .b(new_n21290), .O(new_n21305));
  nor2 g21112(.a(new_n21303), .b(new_n21289), .O(new_n21306));
  nor2 g21113(.a(new_n21306), .b(new_n21305), .O(new_n21307));
  inv1 g21114(.a(new_n21307), .O(new_n21308));
  nor2 g21115(.a(new_n21308), .b(new_n21270), .O(new_n21309));
  nor2 g21116(.a(new_n21307), .b(new_n21269), .O(new_n21310));
  nor2 g21117(.a(new_n21310), .b(new_n21309), .O(new_n21311));
  inv1 g21118(.a(new_n21311), .O(new_n21312));
  nor2 g21119(.a(new_n21159), .b(new_n21155), .O(new_n21313));
  nor2 g21120(.a(new_n21102), .b(new_n21095), .O(new_n21314));
  inv1 g21121(.a(new_n21314), .O(new_n21315));
  nor2 g21122(.a(new_n8476), .b(new_n6274), .O(new_n21316));
  inv1 g21123(.a(new_n21316), .O(new_n21317));
  nor2 g21124(.a(new_n9873), .b(new_n5178), .O(new_n21318));
  nor2 g21125(.a(new_n10320), .b(new_n4954), .O(new_n21319));
  nor2 g21126(.a(new_n21319), .b(new_n21318), .O(new_n21320));
  nor2 g21127(.a(new_n10320), .b(new_n5178), .O(new_n21321));
  inv1 g21128(.a(new_n21321), .O(new_n21322));
  nor2 g21129(.a(new_n21322), .b(new_n21193), .O(new_n21323));
  nor2 g21130(.a(new_n21323), .b(new_n21320), .O(new_n21324));
  nor2 g21131(.a(new_n21324), .b(new_n21317), .O(new_n21325));
  inv1 g21132(.a(new_n21324), .O(new_n21326));
  nor2 g21133(.a(new_n21326), .b(new_n21316), .O(new_n21327));
  nor2 g21134(.a(new_n21327), .b(new_n21325), .O(new_n21328));
  inv1 g21135(.a(new_n21328), .O(new_n21329));
  nor2 g21136(.a(new_n11186), .b(new_n4366), .O(new_n21330));
  nor2 g21137(.a(new_n10468), .b(new_n4682), .O(new_n21331));
  nor2 g21138(.a(new_n21331), .b(new_n21138), .O(new_n21332));
  inv1 g21139(.a(new_n21135), .O(new_n21333));
  nor2 g21140(.a(new_n10895), .b(new_n4682), .O(new_n21334));
  inv1 g21141(.a(new_n21334), .O(new_n21335));
  nor2 g21142(.a(new_n21335), .b(new_n21333), .O(new_n21336));
  nor2 g21143(.a(new_n21336), .b(new_n21332), .O(new_n21337));
  inv1 g21144(.a(new_n21337), .O(new_n21338));
  nor2 g21145(.a(new_n21338), .b(new_n21330), .O(new_n21339));
  inv1 g21146(.a(new_n21330), .O(new_n21340));
  nor2 g21147(.a(new_n21337), .b(new_n21340), .O(new_n21341));
  nor2 g21148(.a(new_n21341), .b(new_n21339), .O(new_n21342));
  nor2 g21149(.a(new_n9156), .b(new_n5796), .O(new_n21343));
  nor2 g21150(.a(new_n21343), .b(new_n20130), .O(new_n21344));
  nor2 g21151(.a(new_n9156), .b(new_n5971), .O(new_n21345));
  inv1 g21152(.a(new_n21345), .O(new_n21346));
  nor2 g21153(.a(new_n21346), .b(new_n21022), .O(new_n21347));
  nor2 g21154(.a(new_n21347), .b(new_n21344), .O(new_n21348));
  nor2 g21155(.a(new_n21348), .b(new_n21170), .O(new_n21349));
  inv1 g21156(.a(new_n21348), .O(new_n21350));
  nor2 g21157(.a(new_n21350), .b(new_n21169), .O(new_n21351));
  nor2 g21158(.a(new_n21351), .b(new_n21349), .O(new_n21352));
  nor2 g21159(.a(new_n21352), .b(new_n21342), .O(new_n21353));
  inv1 g21160(.a(new_n21342), .O(new_n21354));
  inv1 g21161(.a(new_n21352), .O(new_n21355));
  nor2 g21162(.a(new_n21355), .b(new_n21354), .O(new_n21356));
  nor2 g21163(.a(new_n21356), .b(new_n21353), .O(new_n21357));
  nor2 g21164(.a(new_n21357), .b(new_n21329), .O(new_n21358));
  inv1 g21165(.a(new_n21357), .O(new_n21359));
  nor2 g21166(.a(new_n21359), .b(new_n21328), .O(new_n21360));
  nor2 g21167(.a(new_n21360), .b(new_n21358), .O(new_n21361));
  nor2 g21168(.a(new_n21361), .b(new_n21315), .O(new_n21362));
  inv1 g21169(.a(new_n21361), .O(new_n21363));
  nor2 g21170(.a(new_n21363), .b(new_n21314), .O(new_n21364));
  nor2 g21171(.a(new_n21364), .b(new_n21362), .O(new_n21365));
  inv1 g21172(.a(new_n21365), .O(new_n21366));
  nor2 g21173(.a(new_n21151), .b(new_n21120), .O(new_n21367));
  nor2 g21174(.a(new_n21367), .b(new_n21366), .O(new_n21368));
  inv1 g21175(.a(new_n21367), .O(new_n21369));
  nor2 g21176(.a(new_n21369), .b(new_n21365), .O(new_n21370));
  nor2 g21177(.a(new_n21370), .b(new_n21368), .O(new_n21371));
  inv1 g21178(.a(new_n21371), .O(new_n21372));
  nor2 g21179(.a(new_n21372), .b(new_n21313), .O(new_n21373));
  inv1 g21180(.a(new_n21313), .O(new_n21374));
  nor2 g21181(.a(new_n21371), .b(new_n21374), .O(new_n21375));
  nor2 g21182(.a(new_n21375), .b(new_n21373), .O(new_n21376));
  inv1 g21183(.a(new_n21376), .O(new_n21377));
  nor2 g21184(.a(new_n21377), .b(new_n21312), .O(new_n21378));
  nor2 g21185(.a(new_n21376), .b(new_n21311), .O(new_n21379));
  nor2 g21186(.a(new_n21379), .b(new_n21378), .O(new_n21380));
  inv1 g21187(.a(new_n21380), .O(new_n21381));
  nor2 g21188(.a(new_n21381), .b(new_n21240), .O(new_n21382));
  inv1 g21189(.a(new_n21240), .O(new_n21383));
  nor2 g21190(.a(new_n21380), .b(new_n21383), .O(new_n21384));
  nor2 g21191(.a(new_n21384), .b(new_n21382), .O(new_n21385));
  inv1 g21192(.a(new_n21385), .O(new_n21386));
  nor2 g21193(.a(new_n21236), .b(new_n21230), .O(new_n21387));
  nor2 g21194(.a(new_n21387), .b(new_n21386), .O(new_n21388));
  inv1 g21195(.a(new_n21387), .O(new_n21389));
  nor2 g21196(.a(new_n21389), .b(new_n21385), .O(new_n21390));
  nor2 g21197(.a(new_n21390), .b(new_n21388), .O(\asquared[101] ));
  nor2 g21198(.a(new_n21378), .b(new_n21373), .O(new_n21392));
  nor2 g21199(.a(new_n21309), .b(new_n21268), .O(new_n21393));
  nor2 g21200(.a(new_n21262), .b(new_n21253), .O(new_n21394));
  inv1 g21201(.a(new_n21394), .O(new_n21395));
  nor2 g21202(.a(new_n11596), .b(new_n4366), .O(new_n21396));
  nor2 g21203(.a(new_n8946), .b(new_n6274), .O(new_n21397));
  nor2 g21204(.a(new_n8476), .b(new_n6570), .O(new_n21398));
  nor2 g21205(.a(new_n21398), .b(new_n21397), .O(new_n21399));
  nor2 g21206(.a(new_n8946), .b(new_n6570), .O(new_n21400));
  inv1 g21207(.a(new_n21400), .O(new_n21401));
  nor2 g21208(.a(new_n21401), .b(new_n21317), .O(new_n21402));
  nor2 g21209(.a(new_n21402), .b(new_n21399), .O(new_n21403));
  inv1 g21210(.a(new_n21403), .O(new_n21404));
  nor2 g21211(.a(new_n21404), .b(new_n21396), .O(new_n21405));
  inv1 g21212(.a(new_n21396), .O(new_n21406));
  nor2 g21213(.a(new_n21403), .b(new_n21406), .O(new_n21407));
  nor2 g21214(.a(new_n21407), .b(new_n21405), .O(new_n21408));
  nor2 g21215(.a(new_n9873), .b(new_n5393), .O(new_n21409));
  nor2 g21216(.a(new_n21409), .b(new_n21345), .O(new_n21410));
  inv1 g21217(.a(new_n21166), .O(new_n21411));
  nor2 g21218(.a(new_n9873), .b(new_n5971), .O(new_n21412));
  inv1 g21219(.a(new_n21412), .O(new_n21413));
  nor2 g21220(.a(new_n21413), .b(new_n21411), .O(new_n21414));
  nor2 g21221(.a(new_n21414), .b(new_n21410), .O(new_n21415));
  nor2 g21222(.a(new_n21415), .b(new_n21322), .O(new_n21416));
  inv1 g21223(.a(new_n21415), .O(new_n21417));
  nor2 g21224(.a(new_n21417), .b(new_n21321), .O(new_n21418));
  nor2 g21225(.a(new_n21418), .b(new_n21416), .O(new_n21419));
  nor2 g21226(.a(new_n21419), .b(new_n21408), .O(new_n21420));
  inv1 g21227(.a(new_n21408), .O(new_n21421));
  inv1 g21228(.a(new_n21419), .O(new_n21422));
  nor2 g21229(.a(new_n21422), .b(new_n21421), .O(new_n21423));
  nor2 g21230(.a(new_n21423), .b(new_n21420), .O(new_n21424));
  inv1 g21231(.a(new_n21424), .O(new_n21425));
  nor2 g21232(.a(new_n8170), .b(new_n6893), .O(new_n21426));
  inv1 g21233(.a(new_n21426), .O(new_n21427));
  nor2 g21234(.a(new_n9658), .b(new_n5796), .O(new_n21428));
  nor2 g21235(.a(new_n21428), .b(new_n21245), .O(new_n21429));
  nor2 g21236(.a(new_n9658), .b(new_n6958), .O(new_n21430));
  inv1 g21237(.a(new_n21430), .O(new_n21431));
  nor2 g21238(.a(new_n21431), .b(new_n20475), .O(new_n21432));
  nor2 g21239(.a(new_n21432), .b(new_n21429), .O(new_n21433));
  nor2 g21240(.a(new_n21433), .b(new_n21427), .O(new_n21434));
  inv1 g21241(.a(new_n21433), .O(new_n21435));
  nor2 g21242(.a(new_n21435), .b(new_n21426), .O(new_n21436));
  nor2 g21243(.a(new_n21436), .b(new_n21434), .O(new_n21437));
  nor2 g21244(.a(new_n21437), .b(new_n21425), .O(new_n21438));
  inv1 g21245(.a(new_n21437), .O(new_n21439));
  nor2 g21246(.a(new_n21439), .b(new_n21424), .O(new_n21440));
  nor2 g21247(.a(new_n21440), .b(new_n21438), .O(new_n21441));
  nor2 g21248(.a(new_n21441), .b(new_n21395), .O(new_n21442));
  inv1 g21249(.a(new_n21441), .O(new_n21443));
  nor2 g21250(.a(new_n21443), .b(new_n21394), .O(new_n21444));
  nor2 g21251(.a(new_n21444), .b(new_n21442), .O(new_n21445));
  inv1 g21252(.a(new_n21445), .O(new_n21446));
  nor2 g21253(.a(new_n21302), .b(new_n21295), .O(new_n21447));
  nor2 g21254(.a(new_n10468), .b(new_n4954), .O(new_n21448));
  nor2 g21255(.a(new_n21448), .b(new_n21334), .O(new_n21449));
  inv1 g21256(.a(new_n21331), .O(new_n21450));
  nor2 g21257(.a(new_n10895), .b(new_n4954), .O(new_n21451));
  inv1 g21258(.a(new_n21451), .O(new_n21452));
  nor2 g21259(.a(new_n21452), .b(new_n21450), .O(new_n21453));
  nor2 g21260(.a(new_n21453), .b(new_n21449), .O(new_n21454));
  inv1 g21261(.a(new_n21454), .O(new_n21455));
  nor2 g21262(.a(new_n21251), .b(new_n21244), .O(new_n21456));
  inv1 g21263(.a(new_n21456), .O(new_n21457));
  nor2 g21264(.a(new_n21457), .b(new_n21455), .O(new_n21458));
  nor2 g21265(.a(new_n21456), .b(new_n21454), .O(new_n21459));
  nor2 g21266(.a(new_n21459), .b(new_n21458), .O(new_n21460));
  inv1 g21267(.a(new_n21460), .O(new_n21461));
  nor2 g21268(.a(new_n11186), .b(new_n4425), .O(new_n21462));
  inv1 g21269(.a(new_n21462), .O(new_n21463));
  nor2 g21270(.a(new_n7537), .b(\a[50] ), .O(new_n21464));
  nor2 g21271(.a(new_n21464), .b(new_n21463), .O(new_n21465));
  inv1 g21272(.a(new_n21464), .O(new_n21466));
  nor2 g21273(.a(new_n21466), .b(new_n21462), .O(new_n21467));
  nor2 g21274(.a(new_n21467), .b(new_n21465), .O(new_n21468));
  nor2 g21275(.a(new_n21468), .b(new_n21461), .O(new_n21469));
  inv1 g21276(.a(new_n21468), .O(new_n21470));
  nor2 g21277(.a(new_n21470), .b(new_n21460), .O(new_n21471));
  nor2 g21278(.a(new_n21471), .b(new_n21469), .O(new_n21472));
  inv1 g21279(.a(new_n21472), .O(new_n21473));
  nor2 g21280(.a(new_n21473), .b(new_n21447), .O(new_n21474));
  inv1 g21281(.a(new_n21447), .O(new_n21475));
  nor2 g21282(.a(new_n21472), .b(new_n21475), .O(new_n21476));
  nor2 g21283(.a(new_n21476), .b(new_n21474), .O(new_n21477));
  inv1 g21284(.a(new_n21477), .O(new_n21478));
  nor2 g21285(.a(new_n21478), .b(new_n21446), .O(new_n21479));
  nor2 g21286(.a(new_n21477), .b(new_n21445), .O(new_n21480));
  nor2 g21287(.a(new_n21480), .b(new_n21479), .O(new_n21481));
  inv1 g21288(.a(new_n21481), .O(new_n21482));
  nor2 g21289(.a(new_n21482), .b(new_n21393), .O(new_n21483));
  inv1 g21290(.a(new_n21393), .O(new_n21484));
  nor2 g21291(.a(new_n21481), .b(new_n21484), .O(new_n21485));
  nor2 g21292(.a(new_n21485), .b(new_n21483), .O(new_n21486));
  nor2 g21293(.a(new_n21327), .b(new_n21320), .O(new_n21487));
  nor2 g21294(.a(new_n21339), .b(new_n21332), .O(new_n21488));
  nor2 g21295(.a(new_n21488), .b(new_n21487), .O(new_n21489));
  inv1 g21296(.a(new_n21487), .O(new_n21490));
  inv1 g21297(.a(new_n21488), .O(new_n21491));
  nor2 g21298(.a(new_n21491), .b(new_n21490), .O(new_n21492));
  nor2 g21299(.a(new_n21492), .b(new_n21489), .O(new_n21493));
  nor2 g21300(.a(new_n21351), .b(new_n21344), .O(new_n21494));
  nor2 g21301(.a(new_n21494), .b(new_n21493), .O(new_n21495));
  inv1 g21302(.a(new_n21493), .O(new_n21496));
  inv1 g21303(.a(new_n21494), .O(new_n21497));
  nor2 g21304(.a(new_n21497), .b(new_n21496), .O(new_n21498));
  nor2 g21305(.a(new_n21498), .b(new_n21495), .O(new_n21499));
  inv1 g21306(.a(new_n21499), .O(new_n21500));
  nor2 g21307(.a(new_n21282), .b(new_n21276), .O(new_n21501));
  inv1 g21308(.a(new_n21501), .O(new_n21502));
  nor2 g21309(.a(new_n21360), .b(new_n21353), .O(new_n21503));
  inv1 g21310(.a(new_n21503), .O(new_n21504));
  nor2 g21311(.a(new_n21504), .b(new_n21502), .O(new_n21505));
  nor2 g21312(.a(new_n21503), .b(new_n21501), .O(new_n21506));
  nor2 g21313(.a(new_n21506), .b(new_n21505), .O(new_n21507));
  inv1 g21314(.a(new_n21507), .O(new_n21508));
  nor2 g21315(.a(new_n21508), .b(new_n21500), .O(new_n21509));
  nor2 g21316(.a(new_n21507), .b(new_n21499), .O(new_n21510));
  nor2 g21317(.a(new_n21510), .b(new_n21509), .O(new_n21511));
  inv1 g21318(.a(new_n21511), .O(new_n21512));
  nor2 g21319(.a(new_n21368), .b(new_n21364), .O(new_n21513));
  nor2 g21320(.a(new_n21305), .b(new_n21288), .O(new_n21514));
  nor2 g21321(.a(new_n21514), .b(new_n21513), .O(new_n21515));
  inv1 g21322(.a(new_n21513), .O(new_n21516));
  inv1 g21323(.a(new_n21514), .O(new_n21517));
  nor2 g21324(.a(new_n21517), .b(new_n21516), .O(new_n21518));
  nor2 g21325(.a(new_n21518), .b(new_n21515), .O(new_n21519));
  inv1 g21326(.a(new_n21519), .O(new_n21520));
  nor2 g21327(.a(new_n21520), .b(new_n21512), .O(new_n21521));
  nor2 g21328(.a(new_n21519), .b(new_n21511), .O(new_n21522));
  nor2 g21329(.a(new_n21522), .b(new_n21521), .O(new_n21523));
  inv1 g21330(.a(new_n21523), .O(new_n21524));
  nor2 g21331(.a(new_n21524), .b(new_n21486), .O(new_n21525));
  inv1 g21332(.a(new_n21486), .O(new_n21526));
  nor2 g21333(.a(new_n21523), .b(new_n21526), .O(new_n21527));
  nor2 g21334(.a(new_n21527), .b(new_n21525), .O(new_n21528));
  nor2 g21335(.a(new_n21528), .b(new_n21392), .O(new_n21529));
  inv1 g21336(.a(new_n21392), .O(new_n21530));
  inv1 g21337(.a(new_n21528), .O(new_n21531));
  nor2 g21338(.a(new_n21531), .b(new_n21530), .O(new_n21532));
  nor2 g21339(.a(new_n21532), .b(new_n21529), .O(new_n21533));
  inv1 g21340(.a(new_n21533), .O(new_n21534));
  nor2 g21341(.a(new_n21388), .b(new_n21382), .O(new_n21535));
  nor2 g21342(.a(new_n21535), .b(new_n21534), .O(new_n21536));
  inv1 g21343(.a(new_n21535), .O(new_n21537));
  nor2 g21344(.a(new_n21537), .b(new_n21533), .O(new_n21538));
  nor2 g21345(.a(new_n21538), .b(new_n21536), .O(\asquared[102] ));
  nor2 g21346(.a(new_n21467), .b(new_n7537), .O(new_n21540));
  nor2 g21347(.a(new_n21436), .b(new_n21429), .O(new_n21541));
  nor2 g21348(.a(new_n21541), .b(new_n21540), .O(new_n21542));
  inv1 g21349(.a(new_n21540), .O(new_n21543));
  inv1 g21350(.a(new_n21541), .O(new_n21544));
  nor2 g21351(.a(new_n21544), .b(new_n21543), .O(new_n21545));
  nor2 g21352(.a(new_n21545), .b(new_n21542), .O(new_n21546));
  nor2 g21353(.a(new_n21405), .b(new_n21399), .O(new_n21547));
  nor2 g21354(.a(new_n21547), .b(new_n21546), .O(new_n21548));
  inv1 g21355(.a(new_n21546), .O(new_n21549));
  inv1 g21356(.a(new_n21547), .O(new_n21550));
  nor2 g21357(.a(new_n21550), .b(new_n21549), .O(new_n21551));
  nor2 g21358(.a(new_n21551), .b(new_n21548), .O(new_n21552));
  nor2 g21359(.a(new_n21498), .b(new_n21492), .O(new_n21553));
  inv1 g21360(.a(new_n21553), .O(new_n21554));
  nor2 g21361(.a(new_n21554), .b(new_n21552), .O(new_n21555));
  inv1 g21362(.a(new_n21552), .O(new_n21556));
  nor2 g21363(.a(new_n21553), .b(new_n21556), .O(new_n21557));
  nor2 g21364(.a(new_n21557), .b(new_n21555), .O(new_n21558));
  nor2 g21365(.a(new_n21438), .b(new_n21420), .O(new_n21559));
  inv1 g21366(.a(new_n21559), .O(new_n21560));
  nor2 g21367(.a(new_n21560), .b(new_n21558), .O(new_n21561));
  inv1 g21368(.a(new_n21558), .O(new_n21562));
  nor2 g21369(.a(new_n21559), .b(new_n21562), .O(new_n21563));
  nor2 g21370(.a(new_n21563), .b(new_n21561), .O(new_n21564));
  inv1 g21371(.a(new_n21564), .O(new_n21565));
  nor2 g21372(.a(new_n21479), .b(new_n21444), .O(new_n21566));
  nor2 g21373(.a(new_n21509), .b(new_n21506), .O(new_n21567));
  nor2 g21374(.a(new_n21567), .b(new_n21566), .O(new_n21568));
  inv1 g21375(.a(new_n21566), .O(new_n21569));
  inv1 g21376(.a(new_n21567), .O(new_n21570));
  nor2 g21377(.a(new_n21570), .b(new_n21569), .O(new_n21571));
  nor2 g21378(.a(new_n21571), .b(new_n21568), .O(new_n21572));
  inv1 g21379(.a(new_n21572), .O(new_n21573));
  nor2 g21380(.a(new_n21573), .b(new_n21565), .O(new_n21574));
  nor2 g21381(.a(new_n21572), .b(new_n21564), .O(new_n21575));
  nor2 g21382(.a(new_n21575), .b(new_n21574), .O(new_n21576));
  inv1 g21383(.a(new_n21576), .O(new_n21577));
  nor2 g21384(.a(new_n21521), .b(new_n21515), .O(new_n21578));
  nor2 g21385(.a(new_n21474), .b(new_n21469), .O(new_n21579));
  inv1 g21386(.a(new_n21579), .O(new_n21580));
  nor2 g21387(.a(new_n21458), .b(new_n21453), .O(new_n21581));
  inv1 g21388(.a(new_n21581), .O(new_n21582));
  nor2 g21389(.a(new_n21418), .b(new_n21410), .O(new_n21583));
  nor2 g21390(.a(new_n21583), .b(new_n21582), .O(new_n21584));
  inv1 g21391(.a(new_n21583), .O(new_n21585));
  nor2 g21392(.a(new_n21585), .b(new_n21581), .O(new_n21586));
  nor2 g21393(.a(new_n21586), .b(new_n21584), .O(new_n21587));
  inv1 g21394(.a(new_n21587), .O(new_n21588));
  nor2 g21395(.a(new_n11596), .b(new_n4425), .O(new_n21589));
  inv1 g21396(.a(new_n21589), .O(new_n21590));
  nor2 g21397(.a(new_n10468), .b(new_n5178), .O(new_n21591));
  nor2 g21398(.a(new_n21591), .b(new_n21451), .O(new_n21592));
  inv1 g21399(.a(new_n21448), .O(new_n21593));
  nor2 g21400(.a(new_n10895), .b(new_n5178), .O(new_n21594));
  inv1 g21401(.a(new_n21594), .O(new_n21595));
  nor2 g21402(.a(new_n21595), .b(new_n21593), .O(new_n21596));
  nor2 g21403(.a(new_n21596), .b(new_n21592), .O(new_n21597));
  nor2 g21404(.a(new_n21597), .b(new_n21590), .O(new_n21598));
  inv1 g21405(.a(new_n21597), .O(new_n21599));
  nor2 g21406(.a(new_n21599), .b(new_n21589), .O(new_n21600));
  nor2 g21407(.a(new_n21600), .b(new_n21598), .O(new_n21601));
  nor2 g21408(.a(new_n21601), .b(new_n21588), .O(new_n21602));
  inv1 g21409(.a(new_n21601), .O(new_n21603));
  nor2 g21410(.a(new_n21603), .b(new_n21587), .O(new_n21604));
  nor2 g21411(.a(new_n21604), .b(new_n21602), .O(new_n21605));
  nor2 g21412(.a(new_n21605), .b(new_n21580), .O(new_n21606));
  inv1 g21413(.a(new_n21605), .O(new_n21607));
  nor2 g21414(.a(new_n21607), .b(new_n21579), .O(new_n21608));
  nor2 g21415(.a(new_n21608), .b(new_n21606), .O(new_n21609));
  inv1 g21416(.a(new_n21609), .O(new_n21610));
  nor2 g21417(.a(new_n8476), .b(new_n6893), .O(new_n21611));
  inv1 g21418(.a(new_n21611), .O(new_n21612));
  nor2 g21419(.a(new_n8170), .b(new_n6958), .O(new_n21613));
  nor2 g21420(.a(new_n8026), .b(new_n7294), .O(new_n21614));
  nor2 g21421(.a(new_n21614), .b(new_n21613), .O(new_n21615));
  nor2 g21422(.a(new_n8170), .b(new_n7294), .O(new_n21616));
  inv1 g21423(.a(new_n21616), .O(new_n21617));
  nor2 g21424(.a(new_n21617), .b(new_n21246), .O(new_n21618));
  nor2 g21425(.a(new_n21618), .b(new_n21615), .O(new_n21619));
  nor2 g21426(.a(new_n21619), .b(new_n21612), .O(new_n21620));
  inv1 g21427(.a(new_n21619), .O(new_n21621));
  nor2 g21428(.a(new_n21621), .b(new_n21611), .O(new_n21622));
  nor2 g21429(.a(new_n21622), .b(new_n21620), .O(new_n21623));
  inv1 g21430(.a(new_n21623), .O(new_n21624));
  nor2 g21431(.a(new_n9873), .b(new_n5796), .O(new_n21625));
  nor2 g21432(.a(new_n10320), .b(new_n5393), .O(new_n21626));
  nor2 g21433(.a(new_n21626), .b(new_n21625), .O(new_n21627));
  inv1 g21434(.a(new_n21409), .O(new_n21628));
  nor2 g21435(.a(new_n10320), .b(new_n5796), .O(new_n21629));
  inv1 g21436(.a(new_n21629), .O(new_n21630));
  nor2 g21437(.a(new_n21630), .b(new_n21628), .O(new_n21631));
  nor2 g21438(.a(new_n21631), .b(new_n21627), .O(new_n21632));
  inv1 g21439(.a(new_n21632), .O(new_n21633));
  nor2 g21440(.a(new_n21633), .b(new_n16796), .O(new_n21634));
  nor2 g21441(.a(new_n21632), .b(new_n16797), .O(new_n21635));
  nor2 g21442(.a(new_n21635), .b(new_n21634), .O(new_n21636));
  nor2 g21443(.a(new_n9658), .b(new_n5971), .O(new_n21637));
  inv1 g21444(.a(new_n21637), .O(new_n21638));
  nor2 g21445(.a(new_n9156), .b(new_n6274), .O(new_n21639));
  nor2 g21446(.a(new_n21639), .b(new_n21400), .O(new_n21640));
  inv1 g21447(.a(new_n21397), .O(new_n21641));
  nor2 g21448(.a(new_n9156), .b(new_n6570), .O(new_n21642));
  inv1 g21449(.a(new_n21642), .O(new_n21643));
  nor2 g21450(.a(new_n21643), .b(new_n21641), .O(new_n21644));
  nor2 g21451(.a(new_n21644), .b(new_n21640), .O(new_n21645));
  nor2 g21452(.a(new_n21645), .b(new_n21638), .O(new_n21646));
  inv1 g21453(.a(new_n21645), .O(new_n21647));
  nor2 g21454(.a(new_n21647), .b(new_n21637), .O(new_n21648));
  nor2 g21455(.a(new_n21648), .b(new_n21646), .O(new_n21649));
  nor2 g21456(.a(new_n21649), .b(new_n21636), .O(new_n21650));
  inv1 g21457(.a(new_n21636), .O(new_n21651));
  inv1 g21458(.a(new_n21649), .O(new_n21652));
  nor2 g21459(.a(new_n21652), .b(new_n21651), .O(new_n21653));
  nor2 g21460(.a(new_n21653), .b(new_n21650), .O(new_n21654));
  nor2 g21461(.a(new_n21654), .b(new_n21624), .O(new_n21655));
  inv1 g21462(.a(new_n21654), .O(new_n21656));
  nor2 g21463(.a(new_n21656), .b(new_n21623), .O(new_n21657));
  nor2 g21464(.a(new_n21657), .b(new_n21655), .O(new_n21658));
  inv1 g21465(.a(new_n21658), .O(new_n21659));
  nor2 g21466(.a(new_n21659), .b(new_n21610), .O(new_n21660));
  nor2 g21467(.a(new_n21658), .b(new_n21609), .O(new_n21661));
  nor2 g21468(.a(new_n21661), .b(new_n21660), .O(new_n21662));
  inv1 g21469(.a(new_n21662), .O(new_n21663));
  nor2 g21470(.a(new_n21663), .b(new_n21578), .O(new_n21664));
  inv1 g21471(.a(new_n21578), .O(new_n21665));
  nor2 g21472(.a(new_n21662), .b(new_n21665), .O(new_n21666));
  nor2 g21473(.a(new_n21666), .b(new_n21664), .O(new_n21667));
  inv1 g21474(.a(new_n21667), .O(new_n21668));
  nor2 g21475(.a(new_n21668), .b(new_n21577), .O(new_n21669));
  nor2 g21476(.a(new_n21667), .b(new_n21576), .O(new_n21670));
  nor2 g21477(.a(new_n21670), .b(new_n21669), .O(new_n21671));
  nor2 g21478(.a(new_n21527), .b(new_n21485), .O(new_n21672));
  nor2 g21479(.a(new_n21672), .b(new_n21671), .O(new_n21673));
  inv1 g21480(.a(new_n21671), .O(new_n21674));
  inv1 g21481(.a(new_n21672), .O(new_n21675));
  nor2 g21482(.a(new_n21675), .b(new_n21674), .O(new_n21676));
  nor2 g21483(.a(new_n21676), .b(new_n21673), .O(new_n21677));
  inv1 g21484(.a(new_n21677), .O(new_n21678));
  nor2 g21485(.a(new_n21536), .b(new_n21529), .O(new_n21679));
  nor2 g21486(.a(new_n21679), .b(new_n21678), .O(new_n21680));
  inv1 g21487(.a(new_n21679), .O(new_n21681));
  nor2 g21488(.a(new_n21681), .b(new_n21677), .O(new_n21682));
  nor2 g21489(.a(new_n21682), .b(new_n21680), .O(\asquared[103] ));
  nor2 g21490(.a(new_n21669), .b(new_n21664), .O(new_n21684));
  nor2 g21491(.a(new_n21551), .b(new_n21545), .O(new_n21685));
  inv1 g21492(.a(new_n21685), .O(new_n21686));
  nor2 g21493(.a(new_n21602), .b(new_n21586), .O(new_n21687));
  inv1 g21494(.a(new_n21687), .O(new_n21688));
  nor2 g21495(.a(new_n21688), .b(new_n21686), .O(new_n21689));
  nor2 g21496(.a(new_n21687), .b(new_n21685), .O(new_n21690));
  nor2 g21497(.a(new_n21690), .b(new_n21689), .O(new_n21691));
  nor2 g21498(.a(new_n21657), .b(new_n21650), .O(new_n21692));
  inv1 g21499(.a(new_n21692), .O(new_n21693));
  nor2 g21500(.a(new_n21693), .b(new_n21691), .O(new_n21694));
  inv1 g21501(.a(new_n21691), .O(new_n21695));
  nor2 g21502(.a(new_n21692), .b(new_n21695), .O(new_n21696));
  nor2 g21503(.a(new_n21696), .b(new_n21694), .O(new_n21697));
  inv1 g21504(.a(new_n21697), .O(new_n21698));
  nor2 g21505(.a(new_n21660), .b(new_n21608), .O(new_n21699));
  inv1 g21506(.a(new_n21699), .O(new_n21700));
  nor2 g21507(.a(new_n21563), .b(new_n21557), .O(new_n21701));
  inv1 g21508(.a(new_n21701), .O(new_n21702));
  nor2 g21509(.a(new_n21702), .b(new_n21700), .O(new_n21703));
  nor2 g21510(.a(new_n21701), .b(new_n21699), .O(new_n21704));
  nor2 g21511(.a(new_n21704), .b(new_n21703), .O(new_n21705));
  inv1 g21512(.a(new_n21705), .O(new_n21706));
  nor2 g21513(.a(new_n21706), .b(new_n21698), .O(new_n21707));
  nor2 g21514(.a(new_n21705), .b(new_n21697), .O(new_n21708));
  nor2 g21515(.a(new_n21708), .b(new_n21707), .O(new_n21709));
  inv1 g21516(.a(new_n21709), .O(new_n21710));
  nor2 g21517(.a(new_n21574), .b(new_n21568), .O(new_n21711));
  nor2 g21518(.a(new_n11596), .b(new_n4682), .O(new_n21712));
  inv1 g21519(.a(new_n21712), .O(new_n21713));
  nor2 g21520(.a(new_n21622), .b(new_n21615), .O(new_n21714));
  inv1 g21521(.a(new_n21714), .O(new_n21715));
  nor2 g21522(.a(new_n21715), .b(new_n21713), .O(new_n21716));
  nor2 g21523(.a(new_n21714), .b(new_n21712), .O(new_n21717));
  nor2 g21524(.a(new_n21717), .b(new_n21716), .O(new_n21718));
  nor2 g21525(.a(new_n21648), .b(new_n21640), .O(new_n21719));
  nor2 g21526(.a(new_n21719), .b(new_n21718), .O(new_n21720));
  inv1 g21527(.a(new_n21718), .O(new_n21721));
  inv1 g21528(.a(new_n21719), .O(new_n21722));
  nor2 g21529(.a(new_n21722), .b(new_n21721), .O(new_n21723));
  nor2 g21530(.a(new_n21723), .b(new_n21720), .O(new_n21724));
  nor2 g21531(.a(new_n21600), .b(new_n21592), .O(new_n21725));
  nor2 g21532(.a(new_n21634), .b(new_n21627), .O(new_n21726));
  nor2 g21533(.a(new_n21726), .b(new_n21725), .O(new_n21727));
  inv1 g21534(.a(new_n21725), .O(new_n21728));
  inv1 g21535(.a(new_n21726), .O(new_n21729));
  nor2 g21536(.a(new_n21729), .b(new_n21728), .O(new_n21730));
  nor2 g21537(.a(new_n21730), .b(new_n21727), .O(new_n21731));
  inv1 g21538(.a(new_n21731), .O(new_n21732));
  nor2 g21539(.a(new_n21629), .b(new_n21412), .O(new_n21733));
  inv1 g21540(.a(new_n21625), .O(new_n21734));
  nor2 g21541(.a(new_n10320), .b(new_n5971), .O(new_n21735));
  inv1 g21542(.a(new_n21735), .O(new_n21736));
  nor2 g21543(.a(new_n21736), .b(new_n21734), .O(new_n21737));
  nor2 g21544(.a(new_n21737), .b(new_n21733), .O(new_n21738));
  nor2 g21545(.a(new_n21738), .b(new_n21595), .O(new_n21739));
  inv1 g21546(.a(new_n21738), .O(new_n21740));
  nor2 g21547(.a(new_n21740), .b(new_n21594), .O(new_n21741));
  nor2 g21548(.a(new_n21741), .b(new_n21739), .O(new_n21742));
  nor2 g21549(.a(new_n21742), .b(new_n21732), .O(new_n21743));
  inv1 g21550(.a(new_n21742), .O(new_n21744));
  nor2 g21551(.a(new_n21744), .b(new_n21731), .O(new_n21745));
  nor2 g21552(.a(new_n21745), .b(new_n21743), .O(new_n21746));
  nor2 g21553(.a(new_n21746), .b(new_n21724), .O(new_n21747));
  inv1 g21554(.a(new_n21724), .O(new_n21748));
  inv1 g21555(.a(new_n21746), .O(new_n21749));
  nor2 g21556(.a(new_n21749), .b(new_n21748), .O(new_n21750));
  nor2 g21557(.a(new_n21750), .b(new_n21747), .O(new_n21751));
  inv1 g21558(.a(new_n21751), .O(new_n21752));
  nor2 g21559(.a(new_n10468), .b(new_n5393), .O(new_n21753));
  nor2 g21560(.a(new_n9658), .b(new_n6274), .O(new_n21754));
  nor2 g21561(.a(new_n21754), .b(new_n21642), .O(new_n21755));
  inv1 g21562(.a(new_n21639), .O(new_n21756));
  nor2 g21563(.a(new_n9658), .b(new_n6570), .O(new_n21757));
  inv1 g21564(.a(new_n21757), .O(new_n21758));
  nor2 g21565(.a(new_n21758), .b(new_n21756), .O(new_n21759));
  nor2 g21566(.a(new_n21759), .b(new_n21755), .O(new_n21760));
  inv1 g21567(.a(new_n21760), .O(new_n21761));
  nor2 g21568(.a(new_n21761), .b(new_n21753), .O(new_n21762));
  inv1 g21569(.a(new_n21753), .O(new_n21763));
  nor2 g21570(.a(new_n21760), .b(new_n21763), .O(new_n21764));
  nor2 g21571(.a(new_n21764), .b(new_n21762), .O(new_n21765));
  nor2 g21572(.a(new_n8946), .b(new_n6893), .O(new_n21766));
  inv1 g21573(.a(new_n21766), .O(new_n21767));
  nor2 g21574(.a(new_n8476), .b(new_n6958), .O(new_n21768));
  nor2 g21575(.a(new_n21768), .b(new_n21616), .O(new_n21769));
  inv1 g21576(.a(new_n21613), .O(new_n21770));
  nor2 g21577(.a(new_n8476), .b(new_n7294), .O(new_n21771));
  inv1 g21578(.a(new_n21771), .O(new_n21772));
  nor2 g21579(.a(new_n21772), .b(new_n21770), .O(new_n21773));
  nor2 g21580(.a(new_n21773), .b(new_n21769), .O(new_n21774));
  nor2 g21581(.a(new_n21774), .b(new_n21767), .O(new_n21775));
  inv1 g21582(.a(new_n21774), .O(new_n21776));
  nor2 g21583(.a(new_n21776), .b(new_n21766), .O(new_n21777));
  nor2 g21584(.a(new_n21777), .b(new_n21775), .O(new_n21778));
  nor2 g21585(.a(new_n21778), .b(new_n21765), .O(new_n21779));
  inv1 g21586(.a(new_n21765), .O(new_n21780));
  inv1 g21587(.a(new_n21778), .O(new_n21781));
  nor2 g21588(.a(new_n21781), .b(new_n21780), .O(new_n21782));
  nor2 g21589(.a(new_n21782), .b(new_n21779), .O(new_n21783));
  inv1 g21590(.a(new_n21783), .O(new_n21784));
  nor2 g21591(.a(new_n11186), .b(new_n4954), .O(new_n21785));
  inv1 g21592(.a(new_n21785), .O(new_n21786));
  nor2 g21593(.a(new_n8026), .b(\a[51] ), .O(new_n21787));
  nor2 g21594(.a(new_n21787), .b(new_n21786), .O(new_n21788));
  inv1 g21595(.a(new_n21787), .O(new_n21789));
  nor2 g21596(.a(new_n21789), .b(new_n21785), .O(new_n21790));
  nor2 g21597(.a(new_n21790), .b(new_n21788), .O(new_n21791));
  nor2 g21598(.a(new_n21791), .b(new_n21784), .O(new_n21792));
  inv1 g21599(.a(new_n21791), .O(new_n21793));
  nor2 g21600(.a(new_n21793), .b(new_n21783), .O(new_n21794));
  nor2 g21601(.a(new_n21794), .b(new_n21792), .O(new_n21795));
  inv1 g21602(.a(new_n21795), .O(new_n21796));
  nor2 g21603(.a(new_n21796), .b(new_n21752), .O(new_n21797));
  nor2 g21604(.a(new_n21795), .b(new_n21751), .O(new_n21798));
  nor2 g21605(.a(new_n21798), .b(new_n21797), .O(new_n21799));
  inv1 g21606(.a(new_n21799), .O(new_n21800));
  nor2 g21607(.a(new_n21800), .b(new_n21711), .O(new_n21801));
  inv1 g21608(.a(new_n21711), .O(new_n21802));
  nor2 g21609(.a(new_n21799), .b(new_n21802), .O(new_n21803));
  nor2 g21610(.a(new_n21803), .b(new_n21801), .O(new_n21804));
  inv1 g21611(.a(new_n21804), .O(new_n21805));
  nor2 g21612(.a(new_n21805), .b(new_n21710), .O(new_n21806));
  nor2 g21613(.a(new_n21804), .b(new_n21709), .O(new_n21807));
  nor2 g21614(.a(new_n21807), .b(new_n21806), .O(new_n21808));
  inv1 g21615(.a(new_n21808), .O(new_n21809));
  nor2 g21616(.a(new_n21809), .b(new_n21684), .O(new_n21810));
  inv1 g21617(.a(new_n21684), .O(new_n21811));
  nor2 g21618(.a(new_n21808), .b(new_n21811), .O(new_n21812));
  nor2 g21619(.a(new_n21812), .b(new_n21810), .O(new_n21813));
  inv1 g21620(.a(new_n21813), .O(new_n21814));
  nor2 g21621(.a(new_n21680), .b(new_n21676), .O(new_n21815));
  inv1 g21622(.a(new_n21815), .O(new_n21816));
  nor2 g21623(.a(new_n21816), .b(new_n21814), .O(new_n21817));
  nor2 g21624(.a(new_n21815), .b(new_n21813), .O(new_n21818));
  nor2 g21625(.a(new_n21818), .b(new_n21817), .O(new_n21819));
  inv1 g21626(.a(new_n21819), .O(\asquared[104] ));
  nor2 g21627(.a(new_n21806), .b(new_n21801), .O(new_n21821));
  nor2 g21628(.a(new_n21696), .b(new_n21690), .O(new_n21822));
  inv1 g21629(.a(new_n21822), .O(new_n21823));
  nor2 g21630(.a(new_n21797), .b(new_n21750), .O(new_n21824));
  inv1 g21631(.a(new_n21824), .O(new_n21825));
  nor2 g21632(.a(new_n21825), .b(new_n21823), .O(new_n21826));
  nor2 g21633(.a(new_n21824), .b(new_n21822), .O(new_n21827));
  nor2 g21634(.a(new_n21827), .b(new_n21826), .O(new_n21828));
  inv1 g21635(.a(new_n21828), .O(new_n21829));
  nor2 g21636(.a(new_n21723), .b(new_n21716), .O(new_n21830));
  inv1 g21637(.a(new_n21830), .O(new_n21831));
  nor2 g21638(.a(new_n11596), .b(new_n4954), .O(new_n21832));
  nor2 g21639(.a(new_n11186), .b(new_n5178), .O(new_n21833));
  nor2 g21640(.a(new_n21833), .b(new_n21832), .O(new_n21834));
  nor2 g21641(.a(new_n11596), .b(new_n5178), .O(new_n21835));
  inv1 g21642(.a(new_n21835), .O(new_n21836));
  nor2 g21643(.a(new_n21836), .b(new_n21786), .O(new_n21837));
  nor2 g21644(.a(new_n21837), .b(new_n21834), .O(new_n21838));
  inv1 g21645(.a(new_n21838), .O(new_n21839));
  nor2 g21646(.a(new_n21790), .b(new_n8026), .O(new_n21840));
  inv1 g21647(.a(new_n21840), .O(new_n21841));
  nor2 g21648(.a(new_n21841), .b(new_n21839), .O(new_n21842));
  nor2 g21649(.a(new_n21840), .b(new_n21838), .O(new_n21843));
  nor2 g21650(.a(new_n21843), .b(new_n21842), .O(new_n21844));
  nor2 g21651(.a(new_n21844), .b(new_n21831), .O(new_n21845));
  inv1 g21652(.a(new_n21844), .O(new_n21846));
  nor2 g21653(.a(new_n21846), .b(new_n21830), .O(new_n21847));
  nor2 g21654(.a(new_n21847), .b(new_n21845), .O(new_n21848));
  nor2 g21655(.a(new_n21743), .b(new_n21730), .O(new_n21849));
  inv1 g21656(.a(new_n21849), .O(new_n21850));
  nor2 g21657(.a(new_n21850), .b(new_n21848), .O(new_n21851));
  inv1 g21658(.a(new_n21848), .O(new_n21852));
  nor2 g21659(.a(new_n21849), .b(new_n21852), .O(new_n21853));
  nor2 g21660(.a(new_n21853), .b(new_n21851), .O(new_n21854));
  inv1 g21661(.a(new_n21854), .O(new_n21855));
  nor2 g21662(.a(new_n21855), .b(new_n21829), .O(new_n21856));
  nor2 g21663(.a(new_n21854), .b(new_n21828), .O(new_n21857));
  nor2 g21664(.a(new_n21857), .b(new_n21856), .O(new_n21858));
  inv1 g21665(.a(new_n21858), .O(new_n21859));
  nor2 g21666(.a(new_n21707), .b(new_n21704), .O(new_n21860));
  nor2 g21667(.a(new_n21777), .b(new_n21769), .O(new_n21861));
  nor2 g21668(.a(new_n21762), .b(new_n21755), .O(new_n21862));
  nor2 g21669(.a(new_n21862), .b(new_n21861), .O(new_n21863));
  inv1 g21670(.a(new_n21861), .O(new_n21864));
  inv1 g21671(.a(new_n21862), .O(new_n21865));
  nor2 g21672(.a(new_n21865), .b(new_n21864), .O(new_n21866));
  nor2 g21673(.a(new_n21866), .b(new_n21863), .O(new_n21867));
  nor2 g21674(.a(new_n21741), .b(new_n21733), .O(new_n21868));
  nor2 g21675(.a(new_n21868), .b(new_n21867), .O(new_n21869));
  inv1 g21676(.a(new_n21867), .O(new_n21870));
  inv1 g21677(.a(new_n21868), .O(new_n21871));
  nor2 g21678(.a(new_n21871), .b(new_n21870), .O(new_n21872));
  nor2 g21679(.a(new_n21872), .b(new_n21869), .O(new_n21873));
  nor2 g21680(.a(new_n21792), .b(new_n21779), .O(new_n21874));
  inv1 g21681(.a(new_n21874), .O(new_n21875));
  nor2 g21682(.a(new_n21875), .b(new_n21873), .O(new_n21876));
  inv1 g21683(.a(new_n21873), .O(new_n21877));
  nor2 g21684(.a(new_n21874), .b(new_n21877), .O(new_n21878));
  nor2 g21685(.a(new_n21878), .b(new_n21876), .O(new_n21879));
  inv1 g21686(.a(new_n21879), .O(new_n21880));
  nor2 g21687(.a(new_n10468), .b(new_n5796), .O(new_n21881));
  nor2 g21688(.a(new_n10895), .b(new_n5393), .O(new_n21882));
  nor2 g21689(.a(new_n21882), .b(new_n21735), .O(new_n21883));
  inv1 g21690(.a(new_n21626), .O(new_n21884));
  nor2 g21691(.a(new_n10895), .b(new_n5971), .O(new_n21885));
  inv1 g21692(.a(new_n21885), .O(new_n21886));
  nor2 g21693(.a(new_n21886), .b(new_n21884), .O(new_n21887));
  nor2 g21694(.a(new_n21887), .b(new_n21883), .O(new_n21888));
  inv1 g21695(.a(new_n21888), .O(new_n21889));
  nor2 g21696(.a(new_n21889), .b(new_n21881), .O(new_n21890));
  inv1 g21697(.a(new_n21881), .O(new_n21891));
  nor2 g21698(.a(new_n21888), .b(new_n21891), .O(new_n21892));
  nor2 g21699(.a(new_n21892), .b(new_n21890), .O(new_n21893));
  nor2 g21700(.a(new_n9873), .b(new_n6274), .O(new_n21894));
  inv1 g21701(.a(new_n21894), .O(new_n21895));
  nor2 g21702(.a(new_n9156), .b(new_n6893), .O(new_n21896));
  nor2 g21703(.a(new_n21896), .b(new_n21757), .O(new_n21897));
  nor2 g21704(.a(new_n9658), .b(new_n6893), .O(new_n21898));
  inv1 g21705(.a(new_n21898), .O(new_n21899));
  nor2 g21706(.a(new_n21899), .b(new_n21643), .O(new_n21900));
  nor2 g21707(.a(new_n21900), .b(new_n21897), .O(new_n21901));
  nor2 g21708(.a(new_n21901), .b(new_n21895), .O(new_n21902));
  inv1 g21709(.a(new_n21901), .O(new_n21903));
  nor2 g21710(.a(new_n21903), .b(new_n21894), .O(new_n21904));
  nor2 g21711(.a(new_n21904), .b(new_n21902), .O(new_n21905));
  nor2 g21712(.a(new_n21905), .b(new_n21893), .O(new_n21906));
  inv1 g21713(.a(new_n21893), .O(new_n21907));
  inv1 g21714(.a(new_n21905), .O(new_n21908));
  nor2 g21715(.a(new_n21908), .b(new_n21907), .O(new_n21909));
  nor2 g21716(.a(new_n21909), .b(new_n21906), .O(new_n21910));
  inv1 g21717(.a(new_n21910), .O(new_n21911));
  nor2 g21718(.a(new_n8946), .b(new_n6958), .O(new_n21912));
  inv1 g21719(.a(new_n21912), .O(new_n21913));
  nor2 g21720(.a(new_n8170), .b(new_n7537), .O(new_n21914));
  nor2 g21721(.a(new_n21914), .b(new_n21771), .O(new_n21915));
  nor2 g21722(.a(new_n8476), .b(new_n7537), .O(new_n21916));
  inv1 g21723(.a(new_n21916), .O(new_n21917));
  nor2 g21724(.a(new_n21917), .b(new_n21617), .O(new_n21918));
  nor2 g21725(.a(new_n21918), .b(new_n21915), .O(new_n21919));
  nor2 g21726(.a(new_n21919), .b(new_n21913), .O(new_n21920));
  inv1 g21727(.a(new_n21919), .O(new_n21921));
  nor2 g21728(.a(new_n21921), .b(new_n21912), .O(new_n21922));
  nor2 g21729(.a(new_n21922), .b(new_n21920), .O(new_n21923));
  nor2 g21730(.a(new_n21923), .b(new_n21911), .O(new_n21924));
  inv1 g21731(.a(new_n21923), .O(new_n21925));
  nor2 g21732(.a(new_n21925), .b(new_n21910), .O(new_n21926));
  nor2 g21733(.a(new_n21926), .b(new_n21924), .O(new_n21927));
  inv1 g21734(.a(new_n21927), .O(new_n21928));
  nor2 g21735(.a(new_n21928), .b(new_n21880), .O(new_n21929));
  nor2 g21736(.a(new_n21927), .b(new_n21879), .O(new_n21930));
  nor2 g21737(.a(new_n21930), .b(new_n21929), .O(new_n21931));
  inv1 g21738(.a(new_n21931), .O(new_n21932));
  nor2 g21739(.a(new_n21932), .b(new_n21860), .O(new_n21933));
  inv1 g21740(.a(new_n21860), .O(new_n21934));
  nor2 g21741(.a(new_n21931), .b(new_n21934), .O(new_n21935));
  nor2 g21742(.a(new_n21935), .b(new_n21933), .O(new_n21936));
  inv1 g21743(.a(new_n21936), .O(new_n21937));
  nor2 g21744(.a(new_n21937), .b(new_n21859), .O(new_n21938));
  nor2 g21745(.a(new_n21936), .b(new_n21858), .O(new_n21939));
  nor2 g21746(.a(new_n21939), .b(new_n21938), .O(new_n21940));
  inv1 g21747(.a(new_n21940), .O(new_n21941));
  nor2 g21748(.a(new_n21941), .b(new_n21821), .O(new_n21942));
  inv1 g21749(.a(new_n21821), .O(new_n21943));
  nor2 g21750(.a(new_n21940), .b(new_n21943), .O(new_n21944));
  nor2 g21751(.a(new_n21944), .b(new_n21942), .O(new_n21945));
  inv1 g21752(.a(new_n21945), .O(new_n21946));
  nor2 g21753(.a(new_n21815), .b(new_n21812), .O(new_n21947));
  nor2 g21754(.a(new_n21947), .b(new_n21810), .O(new_n21948));
  nor2 g21755(.a(new_n21948), .b(new_n21946), .O(new_n21949));
  inv1 g21756(.a(new_n21948), .O(new_n21950));
  nor2 g21757(.a(new_n21950), .b(new_n21945), .O(new_n21951));
  nor2 g21758(.a(new_n21951), .b(new_n21949), .O(\asquared[105] ));
  nor2 g21759(.a(new_n21904), .b(new_n21897), .O(new_n21953));
  nor2 g21760(.a(new_n21922), .b(new_n21915), .O(new_n21954));
  nor2 g21761(.a(new_n21954), .b(new_n21953), .O(new_n21955));
  inv1 g21762(.a(new_n21953), .O(new_n21956));
  inv1 g21763(.a(new_n21954), .O(new_n21957));
  nor2 g21764(.a(new_n21957), .b(new_n21956), .O(new_n21958));
  nor2 g21765(.a(new_n21958), .b(new_n21955), .O(new_n21959));
  nor2 g21766(.a(new_n21890), .b(new_n21883), .O(new_n21960));
  nor2 g21767(.a(new_n21960), .b(new_n21959), .O(new_n21961));
  inv1 g21768(.a(new_n21959), .O(new_n21962));
  inv1 g21769(.a(new_n21960), .O(new_n21963));
  nor2 g21770(.a(new_n21963), .b(new_n21962), .O(new_n21964));
  nor2 g21771(.a(new_n21964), .b(new_n21961), .O(new_n21965));
  nor2 g21772(.a(new_n21924), .b(new_n21906), .O(new_n21966));
  inv1 g21773(.a(new_n21966), .O(new_n21967));
  nor2 g21774(.a(new_n21967), .b(new_n21965), .O(new_n21968));
  inv1 g21775(.a(new_n21965), .O(new_n21969));
  nor2 g21776(.a(new_n21966), .b(new_n21969), .O(new_n21970));
  nor2 g21777(.a(new_n21970), .b(new_n21968), .O(new_n21971));
  nor2 g21778(.a(new_n21853), .b(new_n21847), .O(new_n21972));
  inv1 g21779(.a(new_n21972), .O(new_n21973));
  nor2 g21780(.a(new_n21973), .b(new_n21971), .O(new_n21974));
  inv1 g21781(.a(new_n21971), .O(new_n21975));
  nor2 g21782(.a(new_n21972), .b(new_n21975), .O(new_n21976));
  nor2 g21783(.a(new_n21976), .b(new_n21974), .O(new_n21977));
  inv1 g21784(.a(new_n21977), .O(new_n21978));
  nor2 g21785(.a(new_n21856), .b(new_n21827), .O(new_n21979));
  nor2 g21786(.a(new_n21979), .b(new_n21978), .O(new_n21980));
  inv1 g21787(.a(new_n21979), .O(new_n21981));
  nor2 g21788(.a(new_n21981), .b(new_n21977), .O(new_n21982));
  nor2 g21789(.a(new_n21982), .b(new_n21980), .O(new_n21983));
  inv1 g21790(.a(new_n21983), .O(new_n21984));
  nor2 g21791(.a(new_n21929), .b(new_n21878), .O(new_n21985));
  nor2 g21792(.a(new_n21872), .b(new_n21866), .O(new_n21986));
  inv1 g21793(.a(new_n21986), .O(new_n21987));
  nor2 g21794(.a(new_n9156), .b(new_n6958), .O(new_n21988));
  inv1 g21795(.a(new_n21988), .O(new_n21989));
  nor2 g21796(.a(new_n8946), .b(new_n7294), .O(new_n21990));
  nor2 g21797(.a(new_n21990), .b(new_n21916), .O(new_n21991));
  nor2 g21798(.a(new_n8946), .b(new_n7537), .O(new_n21992));
  inv1 g21799(.a(new_n21992), .O(new_n21993));
  nor2 g21800(.a(new_n21993), .b(new_n21772), .O(new_n21994));
  nor2 g21801(.a(new_n21994), .b(new_n21991), .O(new_n21995));
  nor2 g21802(.a(new_n21995), .b(new_n21989), .O(new_n21996));
  inv1 g21803(.a(new_n21995), .O(new_n21997));
  nor2 g21804(.a(new_n21997), .b(new_n21988), .O(new_n21998));
  nor2 g21805(.a(new_n21998), .b(new_n21996), .O(new_n21999));
  nor2 g21806(.a(new_n11186), .b(new_n5393), .O(new_n22000));
  inv1 g21807(.a(new_n22000), .O(new_n22001));
  nor2 g21808(.a(new_n8170), .b(\a[52] ), .O(new_n22002));
  nor2 g21809(.a(new_n22002), .b(new_n22001), .O(new_n22003));
  inv1 g21810(.a(new_n22002), .O(new_n22004));
  nor2 g21811(.a(new_n22004), .b(new_n22000), .O(new_n22005));
  nor2 g21812(.a(new_n22005), .b(new_n22003), .O(new_n22006));
  nor2 g21813(.a(new_n22006), .b(new_n21999), .O(new_n22007));
  inv1 g21814(.a(new_n21999), .O(new_n22008));
  inv1 g21815(.a(new_n22006), .O(new_n22009));
  nor2 g21816(.a(new_n22009), .b(new_n22008), .O(new_n22010));
  nor2 g21817(.a(new_n22010), .b(new_n22007), .O(new_n22011));
  nor2 g21818(.a(new_n22011), .b(new_n21987), .O(new_n22012));
  inv1 g21819(.a(new_n22011), .O(new_n22013));
  nor2 g21820(.a(new_n22013), .b(new_n21986), .O(new_n22014));
  nor2 g21821(.a(new_n22014), .b(new_n22012), .O(new_n22015));
  nor2 g21822(.a(new_n10320), .b(new_n6274), .O(new_n22016));
  inv1 g21823(.a(new_n22016), .O(new_n22017));
  nor2 g21824(.a(new_n9873), .b(new_n6570), .O(new_n22018));
  nor2 g21825(.a(new_n22018), .b(new_n21898), .O(new_n22019));
  nor2 g21826(.a(new_n9873), .b(new_n6893), .O(new_n22020));
  inv1 g21827(.a(new_n22020), .O(new_n22021));
  nor2 g21828(.a(new_n22021), .b(new_n21758), .O(new_n22022));
  nor2 g21829(.a(new_n22022), .b(new_n22019), .O(new_n22023));
  nor2 g21830(.a(new_n22023), .b(new_n22017), .O(new_n22024));
  inv1 g21831(.a(new_n22023), .O(new_n22025));
  nor2 g21832(.a(new_n22025), .b(new_n22016), .O(new_n22026));
  nor2 g21833(.a(new_n22026), .b(new_n22024), .O(new_n22027));
  nor2 g21834(.a(new_n10895), .b(new_n5796), .O(new_n22028));
  nor2 g21835(.a(new_n10468), .b(new_n5971), .O(new_n22029));
  nor2 g21836(.a(new_n22029), .b(new_n22028), .O(new_n22030));
  nor2 g21837(.a(new_n21886), .b(new_n21891), .O(new_n22031));
  nor2 g21838(.a(new_n22031), .b(new_n22030), .O(new_n22032));
  nor2 g21839(.a(new_n22032), .b(new_n21836), .O(new_n22033));
  inv1 g21840(.a(new_n22032), .O(new_n22034));
  nor2 g21841(.a(new_n22034), .b(new_n21835), .O(new_n22035));
  nor2 g21842(.a(new_n22035), .b(new_n22033), .O(new_n22036));
  nor2 g21843(.a(new_n21842), .b(new_n21837), .O(new_n22037));
  nor2 g21844(.a(new_n22037), .b(new_n22036), .O(new_n22038));
  inv1 g21845(.a(new_n22036), .O(new_n22039));
  inv1 g21846(.a(new_n22037), .O(new_n22040));
  nor2 g21847(.a(new_n22040), .b(new_n22039), .O(new_n22041));
  nor2 g21848(.a(new_n22041), .b(new_n22038), .O(new_n22042));
  inv1 g21849(.a(new_n22042), .O(new_n22043));
  nor2 g21850(.a(new_n22043), .b(new_n22027), .O(new_n22044));
  inv1 g21851(.a(new_n22027), .O(new_n22045));
  nor2 g21852(.a(new_n22042), .b(new_n22045), .O(new_n22046));
  nor2 g21853(.a(new_n22046), .b(new_n22044), .O(new_n22047));
  nor2 g21854(.a(new_n22047), .b(new_n22015), .O(new_n22048));
  inv1 g21855(.a(new_n22015), .O(new_n22049));
  inv1 g21856(.a(new_n22047), .O(new_n22050));
  nor2 g21857(.a(new_n22050), .b(new_n22049), .O(new_n22051));
  nor2 g21858(.a(new_n22051), .b(new_n22048), .O(new_n22052));
  inv1 g21859(.a(new_n22052), .O(new_n22053));
  nor2 g21860(.a(new_n22053), .b(new_n21985), .O(new_n22054));
  inv1 g21861(.a(new_n21985), .O(new_n22055));
  nor2 g21862(.a(new_n22052), .b(new_n22055), .O(new_n22056));
  nor2 g21863(.a(new_n22056), .b(new_n22054), .O(new_n22057));
  inv1 g21864(.a(new_n22057), .O(new_n22058));
  nor2 g21865(.a(new_n22058), .b(new_n21984), .O(new_n22059));
  nor2 g21866(.a(new_n22057), .b(new_n21983), .O(new_n22060));
  nor2 g21867(.a(new_n22060), .b(new_n22059), .O(new_n22061));
  nor2 g21868(.a(new_n21938), .b(new_n21933), .O(new_n22062));
  inv1 g21869(.a(new_n22062), .O(new_n22063));
  nor2 g21870(.a(new_n22063), .b(new_n22061), .O(new_n22064));
  inv1 g21871(.a(new_n22061), .O(new_n22065));
  nor2 g21872(.a(new_n22062), .b(new_n22065), .O(new_n22066));
  nor2 g21873(.a(new_n22066), .b(new_n22064), .O(new_n22067));
  inv1 g21874(.a(new_n22067), .O(new_n22068));
  nor2 g21875(.a(new_n21949), .b(new_n21942), .O(new_n22069));
  nor2 g21876(.a(new_n22069), .b(new_n22068), .O(new_n22070));
  inv1 g21877(.a(new_n22069), .O(new_n22071));
  nor2 g21878(.a(new_n22071), .b(new_n22067), .O(new_n22072));
  nor2 g21879(.a(new_n22072), .b(new_n22070), .O(\asquared[106] ));
  nor2 g21880(.a(new_n22059), .b(new_n21980), .O(new_n22074));
  nor2 g21881(.a(new_n11596), .b(new_n5393), .O(new_n22075));
  inv1 g21882(.a(new_n22075), .O(new_n22076));
  nor2 g21883(.a(new_n22005), .b(new_n8170), .O(new_n22077));
  inv1 g21884(.a(new_n22077), .O(new_n22078));
  nor2 g21885(.a(new_n22078), .b(new_n22076), .O(new_n22079));
  nor2 g21886(.a(new_n22077), .b(new_n22075), .O(new_n22080));
  nor2 g21887(.a(new_n22080), .b(new_n22079), .O(new_n22081));
  nor2 g21888(.a(new_n21998), .b(new_n21991), .O(new_n22082));
  nor2 g21889(.a(new_n22082), .b(new_n22081), .O(new_n22083));
  inv1 g21890(.a(new_n22081), .O(new_n22084));
  inv1 g21891(.a(new_n22082), .O(new_n22085));
  nor2 g21892(.a(new_n22085), .b(new_n22084), .O(new_n22086));
  nor2 g21893(.a(new_n22086), .b(new_n22083), .O(new_n22087));
  nor2 g21894(.a(new_n22044), .b(new_n22038), .O(new_n22088));
  inv1 g21895(.a(new_n22088), .O(new_n22089));
  nor2 g21896(.a(new_n22089), .b(new_n22087), .O(new_n22090));
  inv1 g21897(.a(new_n22087), .O(new_n22091));
  nor2 g21898(.a(new_n22088), .b(new_n22091), .O(new_n22092));
  nor2 g21899(.a(new_n22092), .b(new_n22090), .O(new_n22093));
  nor2 g21900(.a(new_n22014), .b(new_n22007), .O(new_n22094));
  inv1 g21901(.a(new_n22094), .O(new_n22095));
  nor2 g21902(.a(new_n22095), .b(new_n22093), .O(new_n22096));
  inv1 g21903(.a(new_n22093), .O(new_n22097));
  nor2 g21904(.a(new_n22094), .b(new_n22097), .O(new_n22098));
  nor2 g21905(.a(new_n22098), .b(new_n22096), .O(new_n22099));
  inv1 g21906(.a(new_n22099), .O(new_n22100));
  nor2 g21907(.a(new_n22054), .b(new_n22051), .O(new_n22101));
  nor2 g21908(.a(new_n22101), .b(new_n22100), .O(new_n22102));
  inv1 g21909(.a(new_n22101), .O(new_n22103));
  nor2 g21910(.a(new_n22103), .b(new_n22099), .O(new_n22104));
  nor2 g21911(.a(new_n22104), .b(new_n22102), .O(new_n22105));
  inv1 g21912(.a(new_n22105), .O(new_n22106));
  nor2 g21913(.a(new_n21976), .b(new_n21970), .O(new_n22107));
  nor2 g21914(.a(new_n21964), .b(new_n21958), .O(new_n22108));
  inv1 g21915(.a(new_n22108), .O(new_n22109));
  nor2 g21916(.a(new_n10320), .b(new_n6570), .O(new_n22110));
  nor2 g21917(.a(new_n22020), .b(new_n21430), .O(new_n22111));
  nor2 g21918(.a(new_n9873), .b(new_n6958), .O(new_n22112));
  inv1 g21919(.a(new_n22112), .O(new_n22113));
  nor2 g21920(.a(new_n22113), .b(new_n21899), .O(new_n22114));
  nor2 g21921(.a(new_n22114), .b(new_n22111), .O(new_n22115));
  inv1 g21922(.a(new_n22115), .O(new_n22116));
  nor2 g21923(.a(new_n22116), .b(new_n22110), .O(new_n22117));
  inv1 g21924(.a(new_n22110), .O(new_n22118));
  nor2 g21925(.a(new_n22115), .b(new_n22118), .O(new_n22119));
  nor2 g21926(.a(new_n22119), .b(new_n22117), .O(new_n22120));
  nor2 g21927(.a(new_n9156), .b(new_n7294), .O(new_n22121));
  inv1 g21928(.a(new_n22121), .O(new_n22122));
  nor2 g21929(.a(new_n8476), .b(new_n8026), .O(new_n22123));
  nor2 g21930(.a(new_n22123), .b(new_n21992), .O(new_n22124));
  nor2 g21931(.a(new_n8946), .b(new_n8026), .O(new_n22125));
  inv1 g21932(.a(new_n22125), .O(new_n22126));
  nor2 g21933(.a(new_n22126), .b(new_n21917), .O(new_n22127));
  nor2 g21934(.a(new_n22127), .b(new_n22124), .O(new_n22128));
  nor2 g21935(.a(new_n22128), .b(new_n22122), .O(new_n22129));
  inv1 g21936(.a(new_n22128), .O(new_n22130));
  nor2 g21937(.a(new_n22130), .b(new_n22121), .O(new_n22131));
  nor2 g21938(.a(new_n22131), .b(new_n22129), .O(new_n22132));
  nor2 g21939(.a(new_n22132), .b(new_n22120), .O(new_n22133));
  inv1 g21940(.a(new_n22120), .O(new_n22134));
  inv1 g21941(.a(new_n22132), .O(new_n22135));
  nor2 g21942(.a(new_n22135), .b(new_n22134), .O(new_n22136));
  nor2 g21943(.a(new_n22136), .b(new_n22133), .O(new_n22137));
  nor2 g21944(.a(new_n22137), .b(new_n22109), .O(new_n22138));
  inv1 g21945(.a(new_n22137), .O(new_n22139));
  nor2 g21946(.a(new_n22139), .b(new_n22108), .O(new_n22140));
  nor2 g21947(.a(new_n22140), .b(new_n22138), .O(new_n22141));
  inv1 g21948(.a(new_n22141), .O(new_n22142));
  nor2 g21949(.a(new_n22035), .b(new_n22030), .O(new_n22143));
  nor2 g21950(.a(new_n22026), .b(new_n22019), .O(new_n22144));
  nor2 g21951(.a(new_n22144), .b(new_n22143), .O(new_n22145));
  inv1 g21952(.a(new_n22143), .O(new_n22146));
  inv1 g21953(.a(new_n22144), .O(new_n22147));
  nor2 g21954(.a(new_n22147), .b(new_n22146), .O(new_n22148));
  nor2 g21955(.a(new_n22148), .b(new_n22145), .O(new_n22149));
  inv1 g21956(.a(new_n22149), .O(new_n22150));
  nor2 g21957(.a(new_n11186), .b(new_n5796), .O(new_n22151));
  inv1 g21958(.a(new_n22151), .O(new_n22152));
  nor2 g21959(.a(new_n10468), .b(new_n6274), .O(new_n22153));
  nor2 g21960(.a(new_n22153), .b(new_n21885), .O(new_n22154));
  inv1 g21961(.a(new_n22029), .O(new_n22155));
  nor2 g21962(.a(new_n10895), .b(new_n6274), .O(new_n22156));
  inv1 g21963(.a(new_n22156), .O(new_n22157));
  nor2 g21964(.a(new_n22157), .b(new_n22155), .O(new_n22158));
  nor2 g21965(.a(new_n22158), .b(new_n22154), .O(new_n22159));
  nor2 g21966(.a(new_n22159), .b(new_n22152), .O(new_n22160));
  inv1 g21967(.a(new_n22159), .O(new_n22161));
  nor2 g21968(.a(new_n22161), .b(new_n22151), .O(new_n22162));
  nor2 g21969(.a(new_n22162), .b(new_n22160), .O(new_n22163));
  inv1 g21970(.a(new_n22163), .O(new_n22164));
  nor2 g21971(.a(new_n22164), .b(new_n22150), .O(new_n22165));
  nor2 g21972(.a(new_n22163), .b(new_n22149), .O(new_n22166));
  nor2 g21973(.a(new_n22166), .b(new_n22165), .O(new_n22167));
  nor2 g21974(.a(new_n22167), .b(new_n22142), .O(new_n22168));
  inv1 g21975(.a(new_n22167), .O(new_n22169));
  nor2 g21976(.a(new_n22169), .b(new_n22141), .O(new_n22170));
  nor2 g21977(.a(new_n22170), .b(new_n22168), .O(new_n22171));
  inv1 g21978(.a(new_n22171), .O(new_n22172));
  nor2 g21979(.a(new_n22172), .b(new_n22107), .O(new_n22173));
  inv1 g21980(.a(new_n22107), .O(new_n22174));
  nor2 g21981(.a(new_n22171), .b(new_n22174), .O(new_n22175));
  nor2 g21982(.a(new_n22175), .b(new_n22173), .O(new_n22176));
  inv1 g21983(.a(new_n22176), .O(new_n22177));
  nor2 g21984(.a(new_n22177), .b(new_n22106), .O(new_n22178));
  nor2 g21985(.a(new_n22176), .b(new_n22105), .O(new_n22179));
  nor2 g21986(.a(new_n22179), .b(new_n22178), .O(new_n22180));
  inv1 g21987(.a(new_n22180), .O(new_n22181));
  nor2 g21988(.a(new_n22181), .b(new_n22074), .O(new_n22182));
  inv1 g21989(.a(new_n22074), .O(new_n22183));
  nor2 g21990(.a(new_n22180), .b(new_n22183), .O(new_n22184));
  nor2 g21991(.a(new_n22184), .b(new_n22182), .O(new_n22185));
  inv1 g21992(.a(new_n22185), .O(new_n22186));
  nor2 g21993(.a(new_n22070), .b(new_n22066), .O(new_n22187));
  nor2 g21994(.a(new_n22187), .b(new_n22186), .O(new_n22188));
  inv1 g21995(.a(new_n22187), .O(new_n22189));
  nor2 g21996(.a(new_n22189), .b(new_n22185), .O(new_n22190));
  nor2 g21997(.a(new_n22190), .b(new_n22188), .O(\asquared[107] ));
  nor2 g21998(.a(new_n22178), .b(new_n22102), .O(new_n22192));
  inv1 g21999(.a(new_n22192), .O(new_n22193));
  nor2 g22000(.a(new_n22098), .b(new_n22092), .O(new_n22194));
  inv1 g22001(.a(new_n22194), .O(new_n22195));
  nor2 g22002(.a(new_n10468), .b(new_n6570), .O(new_n22196));
  nor2 g22003(.a(new_n22196), .b(new_n22156), .O(new_n22197));
  inv1 g22004(.a(new_n22153), .O(new_n22198));
  nor2 g22005(.a(new_n10895), .b(new_n6570), .O(new_n22199));
  inv1 g22006(.a(new_n22199), .O(new_n22200));
  nor2 g22007(.a(new_n22200), .b(new_n22198), .O(new_n22201));
  nor2 g22008(.a(new_n22201), .b(new_n22197), .O(new_n22202));
  inv1 g22009(.a(new_n22202), .O(new_n22203));
  nor2 g22010(.a(new_n22131), .b(new_n22124), .O(new_n22204));
  inv1 g22011(.a(new_n22204), .O(new_n22205));
  nor2 g22012(.a(new_n22205), .b(new_n22203), .O(new_n22206));
  nor2 g22013(.a(new_n22204), .b(new_n22202), .O(new_n22207));
  nor2 g22014(.a(new_n22207), .b(new_n22206), .O(new_n22208));
  inv1 g22015(.a(new_n22208), .O(new_n22209));
  nor2 g22016(.a(new_n9658), .b(new_n7294), .O(new_n22210));
  inv1 g22017(.a(new_n22210), .O(new_n22211));
  nor2 g22018(.a(new_n9156), .b(new_n7537), .O(new_n22212));
  nor2 g22019(.a(new_n22212), .b(new_n22125), .O(new_n22213));
  nor2 g22020(.a(new_n9156), .b(new_n8026), .O(new_n22214));
  inv1 g22021(.a(new_n22214), .O(new_n22215));
  nor2 g22022(.a(new_n22215), .b(new_n21993), .O(new_n22216));
  nor2 g22023(.a(new_n22216), .b(new_n22213), .O(new_n22217));
  nor2 g22024(.a(new_n22217), .b(new_n22211), .O(new_n22218));
  inv1 g22025(.a(new_n22217), .O(new_n22219));
  nor2 g22026(.a(new_n22219), .b(new_n22210), .O(new_n22220));
  nor2 g22027(.a(new_n22220), .b(new_n22218), .O(new_n22221));
  nor2 g22028(.a(new_n11186), .b(new_n5971), .O(new_n22222));
  inv1 g22029(.a(new_n22222), .O(new_n22223));
  nor2 g22030(.a(new_n8476), .b(\a[53] ), .O(new_n22224));
  nor2 g22031(.a(new_n22224), .b(new_n22223), .O(new_n22225));
  inv1 g22032(.a(new_n22224), .O(new_n22226));
  nor2 g22033(.a(new_n22226), .b(new_n22222), .O(new_n22227));
  nor2 g22034(.a(new_n22227), .b(new_n22225), .O(new_n22228));
  nor2 g22035(.a(new_n22228), .b(new_n22221), .O(new_n22229));
  inv1 g22036(.a(new_n22221), .O(new_n22230));
  inv1 g22037(.a(new_n22228), .O(new_n22231));
  nor2 g22038(.a(new_n22231), .b(new_n22230), .O(new_n22232));
  nor2 g22039(.a(new_n22232), .b(new_n22229), .O(new_n22233));
  inv1 g22040(.a(new_n22233), .O(new_n22234));
  nor2 g22041(.a(new_n22234), .b(new_n22209), .O(new_n22235));
  nor2 g22042(.a(new_n22233), .b(new_n22208), .O(new_n22236));
  nor2 g22043(.a(new_n22236), .b(new_n22235), .O(new_n22237));
  inv1 g22044(.a(new_n22237), .O(new_n22238));
  nor2 g22045(.a(new_n22162), .b(new_n22154), .O(new_n22239));
  nor2 g22046(.a(new_n22117), .b(new_n22111), .O(new_n22240));
  nor2 g22047(.a(new_n22240), .b(new_n22239), .O(new_n22241));
  inv1 g22048(.a(new_n22239), .O(new_n22242));
  inv1 g22049(.a(new_n22240), .O(new_n22243));
  nor2 g22050(.a(new_n22243), .b(new_n22242), .O(new_n22244));
  nor2 g22051(.a(new_n22244), .b(new_n22241), .O(new_n22245));
  inv1 g22052(.a(new_n22245), .O(new_n22246));
  nor2 g22053(.a(new_n10320), .b(new_n6893), .O(new_n22247));
  inv1 g22054(.a(new_n22247), .O(new_n22248));
  nor2 g22055(.a(new_n11596), .b(new_n5796), .O(new_n22249));
  nor2 g22056(.a(new_n22249), .b(new_n22112), .O(new_n22250));
  nor2 g22057(.a(new_n11596), .b(new_n6958), .O(new_n22251));
  inv1 g22058(.a(new_n22251), .O(new_n22252));
  nor2 g22059(.a(new_n22252), .b(new_n21734), .O(new_n22253));
  nor2 g22060(.a(new_n22253), .b(new_n22250), .O(new_n22254));
  nor2 g22061(.a(new_n22254), .b(new_n22248), .O(new_n22255));
  inv1 g22062(.a(new_n22254), .O(new_n22256));
  nor2 g22063(.a(new_n22256), .b(new_n22247), .O(new_n22257));
  nor2 g22064(.a(new_n22257), .b(new_n22255), .O(new_n22258));
  nor2 g22065(.a(new_n22258), .b(new_n22246), .O(new_n22259));
  inv1 g22066(.a(new_n22258), .O(new_n22260));
  nor2 g22067(.a(new_n22260), .b(new_n22245), .O(new_n22261));
  nor2 g22068(.a(new_n22261), .b(new_n22259), .O(new_n22262));
  inv1 g22069(.a(new_n22262), .O(new_n22263));
  nor2 g22070(.a(new_n22263), .b(new_n22238), .O(new_n22264));
  nor2 g22071(.a(new_n22262), .b(new_n22237), .O(new_n22265));
  nor2 g22072(.a(new_n22265), .b(new_n22264), .O(new_n22266));
  nor2 g22073(.a(new_n22266), .b(new_n22195), .O(new_n22267));
  inv1 g22074(.a(new_n22266), .O(new_n22268));
  nor2 g22075(.a(new_n22268), .b(new_n22194), .O(new_n22269));
  nor2 g22076(.a(new_n22269), .b(new_n22267), .O(new_n22270));
  inv1 g22077(.a(new_n22270), .O(new_n22271));
  nor2 g22078(.a(new_n22173), .b(new_n22168), .O(new_n22272));
  nor2 g22079(.a(new_n22086), .b(new_n22079), .O(new_n22273));
  inv1 g22080(.a(new_n22273), .O(new_n22274));
  nor2 g22081(.a(new_n22165), .b(new_n22145), .O(new_n22275));
  nor2 g22082(.a(new_n22275), .b(new_n22274), .O(new_n22276));
  inv1 g22083(.a(new_n22275), .O(new_n22277));
  nor2 g22084(.a(new_n22277), .b(new_n22273), .O(new_n22278));
  nor2 g22085(.a(new_n22278), .b(new_n22276), .O(new_n22279));
  nor2 g22086(.a(new_n22140), .b(new_n22133), .O(new_n22280));
  inv1 g22087(.a(new_n22280), .O(new_n22281));
  nor2 g22088(.a(new_n22281), .b(new_n22279), .O(new_n22282));
  inv1 g22089(.a(new_n22279), .O(new_n22283));
  nor2 g22090(.a(new_n22280), .b(new_n22283), .O(new_n22284));
  nor2 g22091(.a(new_n22284), .b(new_n22282), .O(new_n22285));
  inv1 g22092(.a(new_n22285), .O(new_n22286));
  nor2 g22093(.a(new_n22286), .b(new_n22272), .O(new_n22287));
  inv1 g22094(.a(new_n22272), .O(new_n22288));
  nor2 g22095(.a(new_n22285), .b(new_n22288), .O(new_n22289));
  nor2 g22096(.a(new_n22289), .b(new_n22287), .O(new_n22290));
  inv1 g22097(.a(new_n22290), .O(new_n22291));
  nor2 g22098(.a(new_n22291), .b(new_n22271), .O(new_n22292));
  nor2 g22099(.a(new_n22290), .b(new_n22270), .O(new_n22293));
  nor2 g22100(.a(new_n22293), .b(new_n22292), .O(new_n22294));
  nor2 g22101(.a(new_n22294), .b(new_n22193), .O(new_n22295));
  inv1 g22102(.a(new_n22294), .O(new_n22296));
  nor2 g22103(.a(new_n22296), .b(new_n22192), .O(new_n22297));
  nor2 g22104(.a(new_n22297), .b(new_n22295), .O(new_n22298));
  inv1 g22105(.a(new_n22298), .O(new_n22299));
  nor2 g22106(.a(new_n22188), .b(new_n22182), .O(new_n22300));
  inv1 g22107(.a(new_n22300), .O(new_n22301));
  nor2 g22108(.a(new_n22301), .b(new_n22299), .O(new_n22302));
  nor2 g22109(.a(new_n22300), .b(new_n22298), .O(new_n22303));
  nor2 g22110(.a(new_n22303), .b(new_n22302), .O(new_n22304));
  inv1 g22111(.a(new_n22304), .O(\asquared[108] ));
  nor2 g22112(.a(new_n22292), .b(new_n22287), .O(new_n22306));
  inv1 g22113(.a(new_n22306), .O(new_n22307));
  nor2 g22114(.a(new_n22269), .b(new_n22264), .O(new_n22308));
  inv1 g22115(.a(new_n22308), .O(new_n22309));
  nor2 g22116(.a(new_n22235), .b(new_n22229), .O(new_n22310));
  nor2 g22117(.a(new_n9658), .b(new_n7537), .O(new_n22311));
  inv1 g22118(.a(new_n22311), .O(new_n22312));
  nor2 g22119(.a(new_n8946), .b(new_n8170), .O(new_n22313));
  nor2 g22120(.a(new_n22313), .b(new_n22214), .O(new_n22314));
  nor2 g22121(.a(new_n9156), .b(new_n8170), .O(new_n22315));
  inv1 g22122(.a(new_n22315), .O(new_n22316));
  nor2 g22123(.a(new_n22316), .b(new_n22126), .O(new_n22317));
  nor2 g22124(.a(new_n22317), .b(new_n22314), .O(new_n22318));
  nor2 g22125(.a(new_n22318), .b(new_n22312), .O(new_n22319));
  inv1 g22126(.a(new_n22318), .O(new_n22320));
  nor2 g22127(.a(new_n22320), .b(new_n22311), .O(new_n22321));
  nor2 g22128(.a(new_n22321), .b(new_n22319), .O(new_n22322));
  nor2 g22129(.a(new_n22259), .b(new_n22244), .O(new_n22323));
  nor2 g22130(.a(new_n22323), .b(new_n22322), .O(new_n22324));
  inv1 g22131(.a(new_n22322), .O(new_n22325));
  inv1 g22132(.a(new_n22323), .O(new_n22326));
  nor2 g22133(.a(new_n22326), .b(new_n22325), .O(new_n22327));
  nor2 g22134(.a(new_n22327), .b(new_n22324), .O(new_n22328));
  inv1 g22135(.a(new_n22328), .O(new_n22329));
  nor2 g22136(.a(new_n22329), .b(new_n22310), .O(new_n22330));
  inv1 g22137(.a(new_n22310), .O(new_n22331));
  nor2 g22138(.a(new_n22328), .b(new_n22331), .O(new_n22332));
  nor2 g22139(.a(new_n22332), .b(new_n22330), .O(new_n22333));
  nor2 g22140(.a(new_n22333), .b(new_n22309), .O(new_n22334));
  inv1 g22141(.a(new_n22333), .O(new_n22335));
  nor2 g22142(.a(new_n22335), .b(new_n22308), .O(new_n22336));
  nor2 g22143(.a(new_n22336), .b(new_n22334), .O(new_n22337));
  inv1 g22144(.a(new_n22337), .O(new_n22338));
  nor2 g22145(.a(new_n22227), .b(new_n8476), .O(new_n22339));
  nor2 g22146(.a(new_n22220), .b(new_n22213), .O(new_n22340));
  nor2 g22147(.a(new_n22340), .b(new_n22339), .O(new_n22341));
  inv1 g22148(.a(new_n22339), .O(new_n22342));
  inv1 g22149(.a(new_n22340), .O(new_n22343));
  nor2 g22150(.a(new_n22343), .b(new_n22342), .O(new_n22344));
  nor2 g22151(.a(new_n22344), .b(new_n22341), .O(new_n22345));
  nor2 g22152(.a(new_n22257), .b(new_n22250), .O(new_n22346));
  nor2 g22153(.a(new_n22346), .b(new_n22345), .O(new_n22347));
  inv1 g22154(.a(new_n22345), .O(new_n22348));
  inv1 g22155(.a(new_n22346), .O(new_n22349));
  nor2 g22156(.a(new_n22349), .b(new_n22348), .O(new_n22350));
  nor2 g22157(.a(new_n22350), .b(new_n22347), .O(new_n22351));
  nor2 g22158(.a(new_n22284), .b(new_n22278), .O(new_n22352));
  inv1 g22159(.a(new_n22352), .O(new_n22353));
  nor2 g22160(.a(new_n22353), .b(new_n22351), .O(new_n22354));
  inv1 g22161(.a(new_n22351), .O(new_n22355));
  nor2 g22162(.a(new_n22352), .b(new_n22355), .O(new_n22356));
  nor2 g22163(.a(new_n22356), .b(new_n22354), .O(new_n22357));
  inv1 g22164(.a(new_n22357), .O(new_n22358));
  nor2 g22165(.a(new_n10468), .b(new_n6893), .O(new_n22359));
  inv1 g22166(.a(new_n22359), .O(new_n22360));
  nor2 g22167(.a(new_n10320), .b(new_n6958), .O(new_n22361));
  nor2 g22168(.a(new_n9873), .b(new_n7294), .O(new_n22362));
  nor2 g22169(.a(new_n22362), .b(new_n22361), .O(new_n22363));
  nor2 g22170(.a(new_n10320), .b(new_n7294), .O(new_n22364));
  inv1 g22171(.a(new_n22364), .O(new_n22365));
  nor2 g22172(.a(new_n22365), .b(new_n22113), .O(new_n22366));
  nor2 g22173(.a(new_n22366), .b(new_n22363), .O(new_n22367));
  nor2 g22174(.a(new_n22367), .b(new_n22360), .O(new_n22368));
  inv1 g22175(.a(new_n22367), .O(new_n22369));
  nor2 g22176(.a(new_n22369), .b(new_n22359), .O(new_n22370));
  nor2 g22177(.a(new_n22370), .b(new_n22368), .O(new_n22371));
  nor2 g22178(.a(new_n11596), .b(new_n5971), .O(new_n22372));
  inv1 g22179(.a(new_n22372), .O(new_n22373));
  nor2 g22180(.a(new_n11186), .b(new_n6274), .O(new_n22374));
  nor2 g22181(.a(new_n22374), .b(new_n22199), .O(new_n22375));
  nor2 g22182(.a(new_n11186), .b(new_n6570), .O(new_n22376));
  inv1 g22183(.a(new_n22376), .O(new_n22377));
  nor2 g22184(.a(new_n22377), .b(new_n22157), .O(new_n22378));
  nor2 g22185(.a(new_n22378), .b(new_n22375), .O(new_n22379));
  nor2 g22186(.a(new_n22379), .b(new_n22373), .O(new_n22380));
  inv1 g22187(.a(new_n22379), .O(new_n22381));
  nor2 g22188(.a(new_n22381), .b(new_n22372), .O(new_n22382));
  nor2 g22189(.a(new_n22382), .b(new_n22380), .O(new_n22383));
  nor2 g22190(.a(new_n22206), .b(new_n22201), .O(new_n22384));
  nor2 g22191(.a(new_n22384), .b(new_n22383), .O(new_n22385));
  inv1 g22192(.a(new_n22383), .O(new_n22386));
  inv1 g22193(.a(new_n22384), .O(new_n22387));
  nor2 g22194(.a(new_n22387), .b(new_n22386), .O(new_n22388));
  nor2 g22195(.a(new_n22388), .b(new_n22385), .O(new_n22389));
  inv1 g22196(.a(new_n22389), .O(new_n22390));
  nor2 g22197(.a(new_n22390), .b(new_n22371), .O(new_n22391));
  inv1 g22198(.a(new_n22371), .O(new_n22392));
  nor2 g22199(.a(new_n22389), .b(new_n22392), .O(new_n22393));
  nor2 g22200(.a(new_n22393), .b(new_n22391), .O(new_n22394));
  inv1 g22201(.a(new_n22394), .O(new_n22395));
  nor2 g22202(.a(new_n22395), .b(new_n22358), .O(new_n22396));
  nor2 g22203(.a(new_n22394), .b(new_n22357), .O(new_n22397));
  nor2 g22204(.a(new_n22397), .b(new_n22396), .O(new_n22398));
  inv1 g22205(.a(new_n22398), .O(new_n22399));
  nor2 g22206(.a(new_n22399), .b(new_n22338), .O(new_n22400));
  nor2 g22207(.a(new_n22398), .b(new_n22337), .O(new_n22401));
  nor2 g22208(.a(new_n22401), .b(new_n22400), .O(new_n22402));
  nor2 g22209(.a(new_n22402), .b(new_n22307), .O(new_n22403));
  inv1 g22210(.a(new_n22402), .O(new_n22404));
  nor2 g22211(.a(new_n22404), .b(new_n22306), .O(new_n22405));
  nor2 g22212(.a(new_n22405), .b(new_n22403), .O(new_n22406));
  inv1 g22213(.a(new_n22406), .O(new_n22407));
  nor2 g22214(.a(new_n22300), .b(new_n22295), .O(new_n22408));
  nor2 g22215(.a(new_n22408), .b(new_n22297), .O(new_n22409));
  nor2 g22216(.a(new_n22409), .b(new_n22407), .O(new_n22410));
  inv1 g22217(.a(new_n22409), .O(new_n22411));
  nor2 g22218(.a(new_n22411), .b(new_n22406), .O(new_n22412));
  nor2 g22219(.a(new_n22412), .b(new_n22410), .O(\asquared[109] ));
  nor2 g22220(.a(new_n22400), .b(new_n22336), .O(new_n22414));
  nor2 g22221(.a(new_n22391), .b(new_n22385), .O(new_n22415));
  inv1 g22222(.a(new_n22415), .O(new_n22416));
  nor2 g22223(.a(new_n22350), .b(new_n22344), .O(new_n22417));
  nor2 g22224(.a(new_n8946), .b(\a[54] ), .O(new_n22418));
  nor2 g22225(.a(new_n22418), .b(new_n22377), .O(new_n22419));
  inv1 g22226(.a(new_n22418), .O(new_n22420));
  nor2 g22227(.a(new_n22420), .b(new_n22376), .O(new_n22421));
  nor2 g22228(.a(new_n22421), .b(new_n22419), .O(new_n22422));
  nor2 g22229(.a(new_n22422), .b(new_n22417), .O(new_n22423));
  inv1 g22230(.a(new_n22417), .O(new_n22424));
  inv1 g22231(.a(new_n22422), .O(new_n22425));
  nor2 g22232(.a(new_n22425), .b(new_n22424), .O(new_n22426));
  nor2 g22233(.a(new_n22426), .b(new_n22423), .O(new_n22427));
  nor2 g22234(.a(new_n22427), .b(new_n22416), .O(new_n22428));
  inv1 g22235(.a(new_n22427), .O(new_n22429));
  nor2 g22236(.a(new_n22429), .b(new_n22415), .O(new_n22430));
  nor2 g22237(.a(new_n22430), .b(new_n22428), .O(new_n22431));
  inv1 g22238(.a(new_n22431), .O(new_n22432));
  nor2 g22239(.a(new_n22396), .b(new_n22356), .O(new_n22433));
  nor2 g22240(.a(new_n22433), .b(new_n22432), .O(new_n22434));
  inv1 g22241(.a(new_n22433), .O(new_n22435));
  nor2 g22242(.a(new_n22435), .b(new_n22431), .O(new_n22436));
  nor2 g22243(.a(new_n22436), .b(new_n22434), .O(new_n22437));
  inv1 g22244(.a(new_n22437), .O(new_n22438));
  nor2 g22245(.a(new_n11596), .b(new_n6274), .O(new_n22439));
  inv1 g22246(.a(new_n22439), .O(new_n22440));
  nor2 g22247(.a(new_n22321), .b(new_n22314), .O(new_n22441));
  inv1 g22248(.a(new_n22441), .O(new_n22442));
  nor2 g22249(.a(new_n22442), .b(new_n22440), .O(new_n22443));
  nor2 g22250(.a(new_n22441), .b(new_n22439), .O(new_n22444));
  nor2 g22251(.a(new_n22444), .b(new_n22443), .O(new_n22445));
  nor2 g22252(.a(new_n22370), .b(new_n22363), .O(new_n22446));
  nor2 g22253(.a(new_n22446), .b(new_n22445), .O(new_n22447));
  inv1 g22254(.a(new_n22445), .O(new_n22448));
  inv1 g22255(.a(new_n22446), .O(new_n22449));
  nor2 g22256(.a(new_n22449), .b(new_n22448), .O(new_n22450));
  nor2 g22257(.a(new_n22450), .b(new_n22447), .O(new_n22451));
  nor2 g22258(.a(new_n22330), .b(new_n22324), .O(new_n22452));
  inv1 g22259(.a(new_n22452), .O(new_n22453));
  nor2 g22260(.a(new_n22453), .b(new_n22451), .O(new_n22454));
  inv1 g22261(.a(new_n22451), .O(new_n22455));
  nor2 g22262(.a(new_n22452), .b(new_n22455), .O(new_n22456));
  nor2 g22263(.a(new_n22456), .b(new_n22454), .O(new_n22457));
  inv1 g22264(.a(new_n22457), .O(new_n22458));
  nor2 g22265(.a(new_n9873), .b(new_n7537), .O(new_n22459));
  inv1 g22266(.a(new_n22459), .O(new_n22460));
  nor2 g22267(.a(new_n9658), .b(new_n8026), .O(new_n22461));
  nor2 g22268(.a(new_n22461), .b(new_n22315), .O(new_n22462));
  nor2 g22269(.a(new_n9658), .b(new_n8170), .O(new_n22463));
  inv1 g22270(.a(new_n22463), .O(new_n22464));
  nor2 g22271(.a(new_n22464), .b(new_n22215), .O(new_n22465));
  nor2 g22272(.a(new_n22465), .b(new_n22462), .O(new_n22466));
  nor2 g22273(.a(new_n22466), .b(new_n22460), .O(new_n22467));
  inv1 g22274(.a(new_n22466), .O(new_n22468));
  nor2 g22275(.a(new_n22468), .b(new_n22459), .O(new_n22469));
  nor2 g22276(.a(new_n22469), .b(new_n22467), .O(new_n22470));
  nor2 g22277(.a(new_n10895), .b(new_n6893), .O(new_n22471));
  inv1 g22278(.a(new_n22471), .O(new_n22472));
  nor2 g22279(.a(new_n10468), .b(new_n6958), .O(new_n22473));
  nor2 g22280(.a(new_n22473), .b(new_n22364), .O(new_n22474));
  inv1 g22281(.a(new_n22361), .O(new_n22475));
  nor2 g22282(.a(new_n10468), .b(new_n7294), .O(new_n22476));
  inv1 g22283(.a(new_n22476), .O(new_n22477));
  nor2 g22284(.a(new_n22477), .b(new_n22475), .O(new_n22478));
  nor2 g22285(.a(new_n22478), .b(new_n22474), .O(new_n22479));
  nor2 g22286(.a(new_n22479), .b(new_n22472), .O(new_n22480));
  inv1 g22287(.a(new_n22479), .O(new_n22481));
  nor2 g22288(.a(new_n22481), .b(new_n22471), .O(new_n22482));
  nor2 g22289(.a(new_n22482), .b(new_n22480), .O(new_n22483));
  nor2 g22290(.a(new_n22382), .b(new_n22375), .O(new_n22484));
  inv1 g22291(.a(new_n22484), .O(new_n22485));
  nor2 g22292(.a(new_n22485), .b(new_n22483), .O(new_n22486));
  inv1 g22293(.a(new_n22483), .O(new_n22487));
  nor2 g22294(.a(new_n22484), .b(new_n22487), .O(new_n22488));
  nor2 g22295(.a(new_n22488), .b(new_n22486), .O(new_n22489));
  inv1 g22296(.a(new_n22489), .O(new_n22490));
  nor2 g22297(.a(new_n22490), .b(new_n22470), .O(new_n22491));
  inv1 g22298(.a(new_n22470), .O(new_n22492));
  nor2 g22299(.a(new_n22489), .b(new_n22492), .O(new_n22493));
  nor2 g22300(.a(new_n22493), .b(new_n22491), .O(new_n22494));
  inv1 g22301(.a(new_n22494), .O(new_n22495));
  nor2 g22302(.a(new_n22495), .b(new_n22458), .O(new_n22496));
  nor2 g22303(.a(new_n22494), .b(new_n22457), .O(new_n22497));
  nor2 g22304(.a(new_n22497), .b(new_n22496), .O(new_n22498));
  inv1 g22305(.a(new_n22498), .O(new_n22499));
  nor2 g22306(.a(new_n22499), .b(new_n22438), .O(new_n22500));
  nor2 g22307(.a(new_n22498), .b(new_n22437), .O(new_n22501));
  nor2 g22308(.a(new_n22501), .b(new_n22500), .O(new_n22502));
  inv1 g22309(.a(new_n22502), .O(new_n22503));
  nor2 g22310(.a(new_n22503), .b(new_n22414), .O(new_n22504));
  inv1 g22311(.a(new_n22414), .O(new_n22505));
  nor2 g22312(.a(new_n22502), .b(new_n22505), .O(new_n22506));
  nor2 g22313(.a(new_n22506), .b(new_n22504), .O(new_n22507));
  inv1 g22314(.a(new_n22507), .O(new_n22508));
  nor2 g22315(.a(new_n22410), .b(new_n22405), .O(new_n22509));
  inv1 g22316(.a(new_n22509), .O(new_n22510));
  nor2 g22317(.a(new_n22510), .b(new_n22508), .O(new_n22511));
  nor2 g22318(.a(new_n22509), .b(new_n22507), .O(new_n22512));
  nor2 g22319(.a(new_n22512), .b(new_n22511), .O(new_n22513));
  inv1 g22320(.a(new_n22513), .O(\asquared[110] ));
  nor2 g22321(.a(new_n22500), .b(new_n22434), .O(new_n22515));
  inv1 g22322(.a(new_n22515), .O(new_n22516));
  nor2 g22323(.a(new_n22491), .b(new_n22486), .O(new_n22517));
  inv1 g22324(.a(new_n22517), .O(new_n22518));
  nor2 g22325(.a(new_n22482), .b(new_n22474), .O(new_n22519));
  nor2 g22326(.a(new_n22469), .b(new_n22462), .O(new_n22520));
  nor2 g22327(.a(new_n22520), .b(new_n22519), .O(new_n22521));
  inv1 g22328(.a(new_n22519), .O(new_n22522));
  inv1 g22329(.a(new_n22520), .O(new_n22523));
  nor2 g22330(.a(new_n22523), .b(new_n22522), .O(new_n22524));
  nor2 g22331(.a(new_n22524), .b(new_n22521), .O(new_n22525));
  inv1 g22332(.a(new_n22525), .O(new_n22526));
  nor2 g22333(.a(new_n10895), .b(new_n6958), .O(new_n22527));
  inv1 g22334(.a(new_n22527), .O(new_n22528));
  nor2 g22335(.a(new_n10320), .b(new_n7537), .O(new_n22529));
  nor2 g22336(.a(new_n22529), .b(new_n22476), .O(new_n22530));
  nor2 g22337(.a(new_n10468), .b(new_n7537), .O(new_n22531));
  inv1 g22338(.a(new_n22531), .O(new_n22532));
  nor2 g22339(.a(new_n22532), .b(new_n22365), .O(new_n22533));
  nor2 g22340(.a(new_n22533), .b(new_n22530), .O(new_n22534));
  nor2 g22341(.a(new_n22534), .b(new_n22528), .O(new_n22535));
  inv1 g22342(.a(new_n22534), .O(new_n22536));
  nor2 g22343(.a(new_n22536), .b(new_n22527), .O(new_n22537));
  nor2 g22344(.a(new_n22537), .b(new_n22535), .O(new_n22538));
  nor2 g22345(.a(new_n22538), .b(new_n22526), .O(new_n22539));
  inv1 g22346(.a(new_n22538), .O(new_n22540));
  nor2 g22347(.a(new_n22540), .b(new_n22525), .O(new_n22541));
  nor2 g22348(.a(new_n22541), .b(new_n22539), .O(new_n22542));
  nor2 g22349(.a(new_n22542), .b(new_n22518), .O(new_n22543));
  inv1 g22350(.a(new_n22542), .O(new_n22544));
  nor2 g22351(.a(new_n22544), .b(new_n22517), .O(new_n22545));
  nor2 g22352(.a(new_n22545), .b(new_n22543), .O(new_n22546));
  nor2 g22353(.a(new_n22430), .b(new_n22423), .O(new_n22547));
  inv1 g22354(.a(new_n22547), .O(new_n22548));
  nor2 g22355(.a(new_n22548), .b(new_n22546), .O(new_n22549));
  inv1 g22356(.a(new_n22546), .O(new_n22550));
  nor2 g22357(.a(new_n22547), .b(new_n22550), .O(new_n22551));
  nor2 g22358(.a(new_n22551), .b(new_n22549), .O(new_n22552));
  inv1 g22359(.a(new_n22552), .O(new_n22553));
  nor2 g22360(.a(new_n22450), .b(new_n22443), .O(new_n22554));
  inv1 g22361(.a(new_n22554), .O(new_n22555));
  nor2 g22362(.a(new_n11186), .b(new_n6893), .O(new_n22556));
  nor2 g22363(.a(new_n11596), .b(new_n6570), .O(new_n22557));
  nor2 g22364(.a(new_n22557), .b(new_n22556), .O(new_n22558));
  nor2 g22365(.a(new_n11596), .b(new_n6893), .O(new_n22559));
  inv1 g22366(.a(new_n22559), .O(new_n22560));
  nor2 g22367(.a(new_n22560), .b(new_n22377), .O(new_n22561));
  nor2 g22368(.a(new_n22561), .b(new_n22558), .O(new_n22562));
  inv1 g22369(.a(new_n22562), .O(new_n22563));
  nor2 g22370(.a(new_n22421), .b(new_n8946), .O(new_n22564));
  inv1 g22371(.a(new_n22564), .O(new_n22565));
  nor2 g22372(.a(new_n22565), .b(new_n22563), .O(new_n22566));
  nor2 g22373(.a(new_n22564), .b(new_n22562), .O(new_n22567));
  nor2 g22374(.a(new_n22567), .b(new_n22566), .O(new_n22568));
  inv1 g22375(.a(new_n22568), .O(new_n22569));
  nor2 g22376(.a(new_n9873), .b(new_n8026), .O(new_n22570));
  inv1 g22377(.a(new_n22570), .O(new_n22571));
  nor2 g22378(.a(new_n9156), .b(new_n8476), .O(new_n22572));
  nor2 g22379(.a(new_n22572), .b(new_n22463), .O(new_n22573));
  nor2 g22380(.a(new_n9658), .b(new_n8476), .O(new_n22574));
  inv1 g22381(.a(new_n22574), .O(new_n22575));
  nor2 g22382(.a(new_n22575), .b(new_n22316), .O(new_n22576));
  nor2 g22383(.a(new_n22576), .b(new_n22573), .O(new_n22577));
  nor2 g22384(.a(new_n22577), .b(new_n22571), .O(new_n22578));
  inv1 g22385(.a(new_n22577), .O(new_n22579));
  nor2 g22386(.a(new_n22579), .b(new_n22570), .O(new_n22580));
  nor2 g22387(.a(new_n22580), .b(new_n22578), .O(new_n22581));
  nor2 g22388(.a(new_n22581), .b(new_n22569), .O(new_n22582));
  inv1 g22389(.a(new_n22581), .O(new_n22583));
  nor2 g22390(.a(new_n22583), .b(new_n22568), .O(new_n22584));
  nor2 g22391(.a(new_n22584), .b(new_n22582), .O(new_n22585));
  nor2 g22392(.a(new_n22585), .b(new_n22555), .O(new_n22586));
  inv1 g22393(.a(new_n22585), .O(new_n22587));
  nor2 g22394(.a(new_n22587), .b(new_n22554), .O(new_n22588));
  nor2 g22395(.a(new_n22588), .b(new_n22586), .O(new_n22589));
  inv1 g22396(.a(new_n22589), .O(new_n22590));
  nor2 g22397(.a(new_n22496), .b(new_n22456), .O(new_n22591));
  nor2 g22398(.a(new_n22591), .b(new_n22590), .O(new_n22592));
  inv1 g22399(.a(new_n22591), .O(new_n22593));
  nor2 g22400(.a(new_n22593), .b(new_n22589), .O(new_n22594));
  nor2 g22401(.a(new_n22594), .b(new_n22592), .O(new_n22595));
  inv1 g22402(.a(new_n22595), .O(new_n22596));
  nor2 g22403(.a(new_n22596), .b(new_n22553), .O(new_n22597));
  nor2 g22404(.a(new_n22595), .b(new_n22552), .O(new_n22598));
  nor2 g22405(.a(new_n22598), .b(new_n22597), .O(new_n22599));
  nor2 g22406(.a(new_n22599), .b(new_n22516), .O(new_n22600));
  inv1 g22407(.a(new_n22599), .O(new_n22601));
  nor2 g22408(.a(new_n22601), .b(new_n22515), .O(new_n22602));
  nor2 g22409(.a(new_n22602), .b(new_n22600), .O(new_n22603));
  inv1 g22410(.a(new_n22603), .O(new_n22604));
  nor2 g22411(.a(new_n22509), .b(new_n22506), .O(new_n22605));
  nor2 g22412(.a(new_n22605), .b(new_n22504), .O(new_n22606));
  nor2 g22413(.a(new_n22606), .b(new_n22604), .O(new_n22607));
  inv1 g22414(.a(new_n22606), .O(new_n22608));
  nor2 g22415(.a(new_n22608), .b(new_n22603), .O(new_n22609));
  nor2 g22416(.a(new_n22609), .b(new_n22607), .O(\asquared[111] ));
  nor2 g22417(.a(new_n22597), .b(new_n22592), .O(new_n22611));
  nor2 g22418(.a(new_n22537), .b(new_n22530), .O(new_n22612));
  nor2 g22419(.a(new_n22580), .b(new_n22573), .O(new_n22613));
  nor2 g22420(.a(new_n22613), .b(new_n22612), .O(new_n22614));
  inv1 g22421(.a(new_n22612), .O(new_n22615));
  inv1 g22422(.a(new_n22613), .O(new_n22616));
  nor2 g22423(.a(new_n22616), .b(new_n22615), .O(new_n22617));
  nor2 g22424(.a(new_n22617), .b(new_n22614), .O(new_n22618));
  nor2 g22425(.a(new_n22566), .b(new_n22561), .O(new_n22619));
  inv1 g22426(.a(new_n22619), .O(new_n22620));
  nor2 g22427(.a(new_n22620), .b(new_n22618), .O(new_n22621));
  inv1 g22428(.a(new_n22618), .O(new_n22622));
  nor2 g22429(.a(new_n22619), .b(new_n22622), .O(new_n22623));
  nor2 g22430(.a(new_n22623), .b(new_n22621), .O(new_n22624));
  nor2 g22431(.a(new_n22539), .b(new_n22524), .O(new_n22625));
  inv1 g22432(.a(new_n22625), .O(new_n22626));
  nor2 g22433(.a(new_n22626), .b(new_n22624), .O(new_n22627));
  inv1 g22434(.a(new_n22624), .O(new_n22628));
  nor2 g22435(.a(new_n22625), .b(new_n22628), .O(new_n22629));
  nor2 g22436(.a(new_n22629), .b(new_n22627), .O(new_n22630));
  nor2 g22437(.a(new_n22588), .b(new_n22582), .O(new_n22631));
  inv1 g22438(.a(new_n22631), .O(new_n22632));
  nor2 g22439(.a(new_n22632), .b(new_n22630), .O(new_n22633));
  inv1 g22440(.a(new_n22630), .O(new_n22634));
  nor2 g22441(.a(new_n22631), .b(new_n22634), .O(new_n22635));
  nor2 g22442(.a(new_n22635), .b(new_n22633), .O(new_n22636));
  inv1 g22443(.a(new_n22636), .O(new_n22637));
  nor2 g22444(.a(new_n22551), .b(new_n22545), .O(new_n22638));
  inv1 g22445(.a(new_n22638), .O(new_n22639));
  nor2 g22446(.a(new_n10320), .b(new_n8026), .O(new_n22640));
  inv1 g22447(.a(new_n22640), .O(new_n22641));
  nor2 g22448(.a(new_n9873), .b(new_n8170), .O(new_n22642));
  nor2 g22449(.a(new_n22642), .b(new_n22574), .O(new_n22643));
  nor2 g22450(.a(new_n9873), .b(new_n8476), .O(new_n22644));
  inv1 g22451(.a(new_n22644), .O(new_n22645));
  nor2 g22452(.a(new_n22645), .b(new_n22464), .O(new_n22646));
  nor2 g22453(.a(new_n22646), .b(new_n22643), .O(new_n22647));
  nor2 g22454(.a(new_n22647), .b(new_n22641), .O(new_n22648));
  inv1 g22455(.a(new_n22647), .O(new_n22649));
  nor2 g22456(.a(new_n22649), .b(new_n22640), .O(new_n22650));
  nor2 g22457(.a(new_n22650), .b(new_n22648), .O(new_n22651));
  inv1 g22458(.a(new_n22651), .O(new_n22652));
  nor2 g22459(.a(new_n10895), .b(new_n7294), .O(new_n22653));
  nor2 g22460(.a(new_n22653), .b(new_n22531), .O(new_n22654));
  nor2 g22461(.a(new_n10895), .b(new_n7537), .O(new_n22655));
  inv1 g22462(.a(new_n22655), .O(new_n22656));
  nor2 g22463(.a(new_n22656), .b(new_n22477), .O(new_n22657));
  nor2 g22464(.a(new_n22657), .b(new_n22654), .O(new_n22658));
  inv1 g22465(.a(new_n22658), .O(new_n22659));
  nor2 g22466(.a(new_n22659), .b(new_n22559), .O(new_n22660));
  nor2 g22467(.a(new_n22658), .b(new_n22560), .O(new_n22661));
  nor2 g22468(.a(new_n22661), .b(new_n22660), .O(new_n22662));
  nor2 g22469(.a(new_n11186), .b(new_n6958), .O(new_n22663));
  inv1 g22470(.a(new_n22663), .O(new_n22664));
  nor2 g22471(.a(new_n9156), .b(\a[55] ), .O(new_n22665));
  nor2 g22472(.a(new_n22665), .b(new_n22664), .O(new_n22666));
  inv1 g22473(.a(new_n22665), .O(new_n22667));
  nor2 g22474(.a(new_n22667), .b(new_n22663), .O(new_n22668));
  nor2 g22475(.a(new_n22668), .b(new_n22666), .O(new_n22669));
  nor2 g22476(.a(new_n22669), .b(new_n22662), .O(new_n22670));
  inv1 g22477(.a(new_n22662), .O(new_n22671));
  inv1 g22478(.a(new_n22669), .O(new_n22672));
  nor2 g22479(.a(new_n22672), .b(new_n22671), .O(new_n22673));
  nor2 g22480(.a(new_n22673), .b(new_n22670), .O(new_n22674));
  nor2 g22481(.a(new_n22674), .b(new_n22652), .O(new_n22675));
  inv1 g22482(.a(new_n22674), .O(new_n22676));
  nor2 g22483(.a(new_n22676), .b(new_n22651), .O(new_n22677));
  nor2 g22484(.a(new_n22677), .b(new_n22675), .O(new_n22678));
  nor2 g22485(.a(new_n22678), .b(new_n22639), .O(new_n22679));
  inv1 g22486(.a(new_n22678), .O(new_n22680));
  nor2 g22487(.a(new_n22680), .b(new_n22638), .O(new_n22681));
  nor2 g22488(.a(new_n22681), .b(new_n22679), .O(new_n22682));
  inv1 g22489(.a(new_n22682), .O(new_n22683));
  nor2 g22490(.a(new_n22683), .b(new_n22637), .O(new_n22684));
  nor2 g22491(.a(new_n22682), .b(new_n22636), .O(new_n22685));
  nor2 g22492(.a(new_n22685), .b(new_n22684), .O(new_n22686));
  inv1 g22493(.a(new_n22686), .O(new_n22687));
  nor2 g22494(.a(new_n22687), .b(new_n22611), .O(new_n22688));
  inv1 g22495(.a(new_n22611), .O(new_n22689));
  nor2 g22496(.a(new_n22686), .b(new_n22689), .O(new_n22690));
  nor2 g22497(.a(new_n22690), .b(new_n22688), .O(new_n22691));
  inv1 g22498(.a(new_n22691), .O(new_n22692));
  nor2 g22499(.a(new_n22607), .b(new_n22602), .O(new_n22693));
  inv1 g22500(.a(new_n22693), .O(new_n22694));
  nor2 g22501(.a(new_n22694), .b(new_n22692), .O(new_n22695));
  nor2 g22502(.a(new_n22693), .b(new_n22691), .O(new_n22696));
  nor2 g22503(.a(new_n22696), .b(new_n22695), .O(new_n22697));
  inv1 g22504(.a(new_n22697), .O(\asquared[112] ));
  nor2 g22505(.a(new_n22684), .b(new_n22681), .O(new_n22699));
  inv1 g22506(.a(new_n22699), .O(new_n22700));
  nor2 g22507(.a(new_n22635), .b(new_n22629), .O(new_n22701));
  inv1 g22508(.a(new_n22701), .O(new_n22702));
  nor2 g22509(.a(new_n10320), .b(new_n8170), .O(new_n22703));
  inv1 g22510(.a(new_n22703), .O(new_n22704));
  nor2 g22511(.a(new_n9658), .b(new_n8946), .O(new_n22705));
  nor2 g22512(.a(new_n22705), .b(new_n22644), .O(new_n22706));
  nor2 g22513(.a(new_n9873), .b(new_n8946), .O(new_n22707));
  inv1 g22514(.a(new_n22707), .O(new_n22708));
  nor2 g22515(.a(new_n22708), .b(new_n22575), .O(new_n22709));
  nor2 g22516(.a(new_n22709), .b(new_n22706), .O(new_n22710));
  nor2 g22517(.a(new_n22710), .b(new_n22704), .O(new_n22711));
  inv1 g22518(.a(new_n22710), .O(new_n22712));
  nor2 g22519(.a(new_n22712), .b(new_n22703), .O(new_n22713));
  nor2 g22520(.a(new_n22713), .b(new_n22711), .O(new_n22714));
  nor2 g22521(.a(new_n10468), .b(new_n8026), .O(new_n22715));
  nor2 g22522(.a(new_n22715), .b(new_n22655), .O(new_n22716));
  nor2 g22523(.a(new_n10895), .b(new_n8026), .O(new_n22717));
  inv1 g22524(.a(new_n22717), .O(new_n22718));
  nor2 g22525(.a(new_n22718), .b(new_n22532), .O(new_n22719));
  nor2 g22526(.a(new_n22719), .b(new_n22716), .O(new_n22720));
  nor2 g22527(.a(new_n22720), .b(new_n22252), .O(new_n22721));
  inv1 g22528(.a(new_n22720), .O(new_n22722));
  nor2 g22529(.a(new_n22722), .b(new_n22251), .O(new_n22723));
  nor2 g22530(.a(new_n22723), .b(new_n22721), .O(new_n22724));
  nor2 g22531(.a(new_n22660), .b(new_n22654), .O(new_n22725));
  inv1 g22532(.a(new_n22725), .O(new_n22726));
  nor2 g22533(.a(new_n22726), .b(new_n22724), .O(new_n22727));
  inv1 g22534(.a(new_n22724), .O(new_n22728));
  nor2 g22535(.a(new_n22725), .b(new_n22728), .O(new_n22729));
  nor2 g22536(.a(new_n22729), .b(new_n22727), .O(new_n22730));
  inv1 g22537(.a(new_n22730), .O(new_n22731));
  nor2 g22538(.a(new_n22731), .b(new_n22714), .O(new_n22732));
  inv1 g22539(.a(new_n22714), .O(new_n22733));
  nor2 g22540(.a(new_n22730), .b(new_n22733), .O(new_n22734));
  nor2 g22541(.a(new_n22734), .b(new_n22732), .O(new_n22735));
  nor2 g22542(.a(new_n22735), .b(new_n22702), .O(new_n22736));
  inv1 g22543(.a(new_n22735), .O(new_n22737));
  nor2 g22544(.a(new_n22737), .b(new_n22701), .O(new_n22738));
  nor2 g22545(.a(new_n22738), .b(new_n22736), .O(new_n22739));
  inv1 g22546(.a(new_n22739), .O(new_n22740));
  nor2 g22547(.a(new_n11186), .b(new_n7294), .O(new_n22741));
  inv1 g22548(.a(new_n22741), .O(new_n22742));
  nor2 g22549(.a(new_n22668), .b(new_n9156), .O(new_n22743));
  inv1 g22550(.a(new_n22743), .O(new_n22744));
  nor2 g22551(.a(new_n22744), .b(new_n22742), .O(new_n22745));
  nor2 g22552(.a(new_n22743), .b(new_n22741), .O(new_n22746));
  nor2 g22553(.a(new_n22746), .b(new_n22745), .O(new_n22747));
  nor2 g22554(.a(new_n22650), .b(new_n22643), .O(new_n22748));
  nor2 g22555(.a(new_n22748), .b(new_n22747), .O(new_n22749));
  inv1 g22556(.a(new_n22747), .O(new_n22750));
  inv1 g22557(.a(new_n22748), .O(new_n22751));
  nor2 g22558(.a(new_n22751), .b(new_n22750), .O(new_n22752));
  nor2 g22559(.a(new_n22752), .b(new_n22749), .O(new_n22753));
  inv1 g22560(.a(new_n22753), .O(new_n22754));
  nor2 g22561(.a(new_n22623), .b(new_n22617), .O(new_n22755));
  inv1 g22562(.a(new_n22755), .O(new_n22756));
  nor2 g22563(.a(new_n22677), .b(new_n22670), .O(new_n22757));
  inv1 g22564(.a(new_n22757), .O(new_n22758));
  nor2 g22565(.a(new_n22758), .b(new_n22756), .O(new_n22759));
  nor2 g22566(.a(new_n22757), .b(new_n22755), .O(new_n22760));
  nor2 g22567(.a(new_n22760), .b(new_n22759), .O(new_n22761));
  inv1 g22568(.a(new_n22761), .O(new_n22762));
  nor2 g22569(.a(new_n22762), .b(new_n22754), .O(new_n22763));
  nor2 g22570(.a(new_n22761), .b(new_n22753), .O(new_n22764));
  nor2 g22571(.a(new_n22764), .b(new_n22763), .O(new_n22765));
  inv1 g22572(.a(new_n22765), .O(new_n22766));
  nor2 g22573(.a(new_n22766), .b(new_n22740), .O(new_n22767));
  nor2 g22574(.a(new_n22765), .b(new_n22739), .O(new_n22768));
  nor2 g22575(.a(new_n22768), .b(new_n22767), .O(new_n22769));
  nor2 g22576(.a(new_n22769), .b(new_n22700), .O(new_n22770));
  inv1 g22577(.a(new_n22769), .O(new_n22771));
  nor2 g22578(.a(new_n22771), .b(new_n22699), .O(new_n22772));
  nor2 g22579(.a(new_n22772), .b(new_n22770), .O(new_n22773));
  inv1 g22580(.a(new_n22773), .O(new_n22774));
  nor2 g22581(.a(new_n22693), .b(new_n22690), .O(new_n22775));
  nor2 g22582(.a(new_n22775), .b(new_n22688), .O(new_n22776));
  nor2 g22583(.a(new_n22776), .b(new_n22774), .O(new_n22777));
  inv1 g22584(.a(new_n22776), .O(new_n22778));
  nor2 g22585(.a(new_n22778), .b(new_n22773), .O(new_n22779));
  nor2 g22586(.a(new_n22779), .b(new_n22777), .O(\asquared[113] ));
  nor2 g22587(.a(new_n22767), .b(new_n22738), .O(new_n22781));
  inv1 g22588(.a(new_n22781), .O(new_n22782));
  nor2 g22589(.a(new_n22752), .b(new_n22745), .O(new_n22783));
  inv1 g22590(.a(new_n22783), .O(new_n22784));
  nor2 g22591(.a(new_n10468), .b(new_n8170), .O(new_n22785));
  nor2 g22592(.a(new_n22785), .b(new_n22717), .O(new_n22786));
  inv1 g22593(.a(new_n22715), .O(new_n22787));
  nor2 g22594(.a(new_n10895), .b(new_n8170), .O(new_n22788));
  inv1 g22595(.a(new_n22788), .O(new_n22789));
  nor2 g22596(.a(new_n22789), .b(new_n22787), .O(new_n22790));
  nor2 g22597(.a(new_n22790), .b(new_n22786), .O(new_n22791));
  inv1 g22598(.a(new_n22791), .O(new_n22792));
  nor2 g22599(.a(new_n22713), .b(new_n22706), .O(new_n22793));
  inv1 g22600(.a(new_n22793), .O(new_n22794));
  nor2 g22601(.a(new_n22794), .b(new_n22792), .O(new_n22795));
  nor2 g22602(.a(new_n22793), .b(new_n22791), .O(new_n22796));
  nor2 g22603(.a(new_n22796), .b(new_n22795), .O(new_n22797));
  nor2 g22604(.a(new_n22797), .b(new_n22784), .O(new_n22798));
  inv1 g22605(.a(new_n22797), .O(new_n22799));
  nor2 g22606(.a(new_n22799), .b(new_n22783), .O(new_n22800));
  nor2 g22607(.a(new_n22800), .b(new_n22798), .O(new_n22801));
  nor2 g22608(.a(new_n22732), .b(new_n22727), .O(new_n22802));
  inv1 g22609(.a(new_n22802), .O(new_n22803));
  nor2 g22610(.a(new_n22803), .b(new_n22801), .O(new_n22804));
  inv1 g22611(.a(new_n22801), .O(new_n22805));
  nor2 g22612(.a(new_n22802), .b(new_n22805), .O(new_n22806));
  nor2 g22613(.a(new_n22806), .b(new_n22804), .O(new_n22807));
  nor2 g22614(.a(new_n22763), .b(new_n22760), .O(new_n22808));
  nor2 g22615(.a(new_n11596), .b(new_n7294), .O(new_n22809));
  inv1 g22616(.a(new_n22809), .O(new_n22810));
  nor2 g22617(.a(new_n10320), .b(new_n8476), .O(new_n22811));
  nor2 g22618(.a(new_n22811), .b(new_n22707), .O(new_n22812));
  nor2 g22619(.a(new_n10320), .b(new_n8946), .O(new_n22813));
  inv1 g22620(.a(new_n22813), .O(new_n22814));
  nor2 g22621(.a(new_n22814), .b(new_n22645), .O(new_n22815));
  nor2 g22622(.a(new_n22815), .b(new_n22812), .O(new_n22816));
  nor2 g22623(.a(new_n22816), .b(new_n22810), .O(new_n22817));
  inv1 g22624(.a(new_n22816), .O(new_n22818));
  nor2 g22625(.a(new_n22818), .b(new_n22809), .O(new_n22819));
  nor2 g22626(.a(new_n22819), .b(new_n22817), .O(new_n22820));
  nor2 g22627(.a(new_n22723), .b(new_n22716), .O(new_n22821));
  inv1 g22628(.a(new_n22821), .O(new_n22822));
  nor2 g22629(.a(new_n22822), .b(new_n22820), .O(new_n22823));
  inv1 g22630(.a(new_n22820), .O(new_n22824));
  nor2 g22631(.a(new_n22821), .b(new_n22824), .O(new_n22825));
  nor2 g22632(.a(new_n22825), .b(new_n22823), .O(new_n22826));
  inv1 g22633(.a(new_n22826), .O(new_n22827));
  nor2 g22634(.a(new_n11186), .b(new_n7537), .O(new_n22828));
  inv1 g22635(.a(new_n22828), .O(new_n22829));
  nor2 g22636(.a(new_n9658), .b(\a[56] ), .O(new_n22830));
  nor2 g22637(.a(new_n22830), .b(new_n22829), .O(new_n22831));
  inv1 g22638(.a(new_n22830), .O(new_n22832));
  nor2 g22639(.a(new_n22832), .b(new_n22828), .O(new_n22833));
  nor2 g22640(.a(new_n22833), .b(new_n22831), .O(new_n22834));
  nor2 g22641(.a(new_n22834), .b(new_n22827), .O(new_n22835));
  inv1 g22642(.a(new_n22834), .O(new_n22836));
  nor2 g22643(.a(new_n22836), .b(new_n22826), .O(new_n22837));
  nor2 g22644(.a(new_n22837), .b(new_n22835), .O(new_n22838));
  inv1 g22645(.a(new_n22838), .O(new_n22839));
  nor2 g22646(.a(new_n22839), .b(new_n22808), .O(new_n22840));
  inv1 g22647(.a(new_n22808), .O(new_n22841));
  nor2 g22648(.a(new_n22838), .b(new_n22841), .O(new_n22842));
  nor2 g22649(.a(new_n22842), .b(new_n22840), .O(new_n22843));
  nor2 g22650(.a(new_n22843), .b(new_n22807), .O(new_n22844));
  inv1 g22651(.a(new_n22807), .O(new_n22845));
  inv1 g22652(.a(new_n22843), .O(new_n22846));
  nor2 g22653(.a(new_n22846), .b(new_n22845), .O(new_n22847));
  nor2 g22654(.a(new_n22847), .b(new_n22844), .O(new_n22848));
  nor2 g22655(.a(new_n22848), .b(new_n22782), .O(new_n22849));
  inv1 g22656(.a(new_n22848), .O(new_n22850));
  nor2 g22657(.a(new_n22850), .b(new_n22781), .O(new_n22851));
  nor2 g22658(.a(new_n22851), .b(new_n22849), .O(new_n22852));
  inv1 g22659(.a(new_n22852), .O(new_n22853));
  nor2 g22660(.a(new_n22777), .b(new_n22772), .O(new_n22854));
  inv1 g22661(.a(new_n22854), .O(new_n22855));
  nor2 g22662(.a(new_n22855), .b(new_n22853), .O(new_n22856));
  nor2 g22663(.a(new_n22854), .b(new_n22852), .O(new_n22857));
  nor2 g22664(.a(new_n22857), .b(new_n22856), .O(new_n22858));
  inv1 g22665(.a(new_n22858), .O(\asquared[114] ));
  nor2 g22666(.a(new_n22847), .b(new_n22840), .O(new_n22860));
  inv1 g22667(.a(new_n22860), .O(new_n22861));
  nor2 g22668(.a(new_n22833), .b(new_n9658), .O(new_n22862));
  nor2 g22669(.a(new_n22819), .b(new_n22812), .O(new_n22863));
  nor2 g22670(.a(new_n22863), .b(new_n22862), .O(new_n22864));
  inv1 g22671(.a(new_n22862), .O(new_n22865));
  inv1 g22672(.a(new_n22863), .O(new_n22866));
  nor2 g22673(.a(new_n22866), .b(new_n22865), .O(new_n22867));
  nor2 g22674(.a(new_n22867), .b(new_n22864), .O(new_n22868));
  nor2 g22675(.a(new_n22795), .b(new_n22790), .O(new_n22869));
  inv1 g22676(.a(new_n22869), .O(new_n22870));
  nor2 g22677(.a(new_n22870), .b(new_n22868), .O(new_n22871));
  inv1 g22678(.a(new_n22868), .O(new_n22872));
  nor2 g22679(.a(new_n22869), .b(new_n22872), .O(new_n22873));
  nor2 g22680(.a(new_n22873), .b(new_n22871), .O(new_n22874));
  nor2 g22681(.a(new_n22806), .b(new_n22800), .O(new_n22875));
  inv1 g22682(.a(new_n22875), .O(new_n22876));
  nor2 g22683(.a(new_n22876), .b(new_n22874), .O(new_n22877));
  inv1 g22684(.a(new_n22874), .O(new_n22878));
  nor2 g22685(.a(new_n22875), .b(new_n22878), .O(new_n22879));
  nor2 g22686(.a(new_n22879), .b(new_n22877), .O(new_n22880));
  inv1 g22687(.a(new_n22880), .O(new_n22881));
  nor2 g22688(.a(new_n22835), .b(new_n22823), .O(new_n22882));
  inv1 g22689(.a(new_n22882), .O(new_n22883));
  nor2 g22690(.a(new_n11596), .b(new_n7537), .O(new_n22884));
  nor2 g22691(.a(new_n11186), .b(new_n8026), .O(new_n22885));
  nor2 g22692(.a(new_n22885), .b(new_n22788), .O(new_n22886));
  nor2 g22693(.a(new_n11186), .b(new_n8170), .O(new_n22887));
  inv1 g22694(.a(new_n22887), .O(new_n22888));
  nor2 g22695(.a(new_n22888), .b(new_n22718), .O(new_n22889));
  nor2 g22696(.a(new_n22889), .b(new_n22886), .O(new_n22890));
  inv1 g22697(.a(new_n22890), .O(new_n22891));
  nor2 g22698(.a(new_n22891), .b(new_n22884), .O(new_n22892));
  inv1 g22699(.a(new_n22884), .O(new_n22893));
  nor2 g22700(.a(new_n22890), .b(new_n22893), .O(new_n22894));
  nor2 g22701(.a(new_n22894), .b(new_n22892), .O(new_n22895));
  nor2 g22702(.a(new_n10468), .b(new_n8476), .O(new_n22896));
  inv1 g22703(.a(new_n22896), .O(new_n22897));
  nor2 g22704(.a(new_n9873), .b(new_n9156), .O(new_n22898));
  nor2 g22705(.a(new_n22898), .b(new_n22813), .O(new_n22899));
  nor2 g22706(.a(new_n10320), .b(new_n9156), .O(new_n22900));
  inv1 g22707(.a(new_n22900), .O(new_n22901));
  nor2 g22708(.a(new_n22901), .b(new_n22708), .O(new_n22902));
  nor2 g22709(.a(new_n22902), .b(new_n22899), .O(new_n22903));
  nor2 g22710(.a(new_n22903), .b(new_n22897), .O(new_n22904));
  inv1 g22711(.a(new_n22903), .O(new_n22905));
  nor2 g22712(.a(new_n22905), .b(new_n22896), .O(new_n22906));
  nor2 g22713(.a(new_n22906), .b(new_n22904), .O(new_n22907));
  nor2 g22714(.a(new_n22907), .b(new_n22895), .O(new_n22908));
  inv1 g22715(.a(new_n22895), .O(new_n22909));
  inv1 g22716(.a(new_n22907), .O(new_n22910));
  nor2 g22717(.a(new_n22910), .b(new_n22909), .O(new_n22911));
  nor2 g22718(.a(new_n22911), .b(new_n22908), .O(new_n22912));
  nor2 g22719(.a(new_n22912), .b(new_n22883), .O(new_n22913));
  inv1 g22720(.a(new_n22912), .O(new_n22914));
  nor2 g22721(.a(new_n22914), .b(new_n22882), .O(new_n22915));
  nor2 g22722(.a(new_n22915), .b(new_n22913), .O(new_n22916));
  inv1 g22723(.a(new_n22916), .O(new_n22917));
  nor2 g22724(.a(new_n22917), .b(new_n22881), .O(new_n22918));
  nor2 g22725(.a(new_n22916), .b(new_n22880), .O(new_n22919));
  nor2 g22726(.a(new_n22919), .b(new_n22918), .O(new_n22920));
  nor2 g22727(.a(new_n22920), .b(new_n22861), .O(new_n22921));
  inv1 g22728(.a(new_n22920), .O(new_n22922));
  nor2 g22729(.a(new_n22922), .b(new_n22860), .O(new_n22923));
  nor2 g22730(.a(new_n22923), .b(new_n22921), .O(new_n22924));
  inv1 g22731(.a(new_n22924), .O(new_n22925));
  nor2 g22732(.a(new_n22854), .b(new_n22849), .O(new_n22926));
  nor2 g22733(.a(new_n22926), .b(new_n22851), .O(new_n22927));
  nor2 g22734(.a(new_n22927), .b(new_n22925), .O(new_n22928));
  inv1 g22735(.a(new_n22927), .O(new_n22929));
  nor2 g22736(.a(new_n22929), .b(new_n22924), .O(new_n22930));
  nor2 g22737(.a(new_n22930), .b(new_n22928), .O(\asquared[115] ));
  nor2 g22738(.a(new_n22918), .b(new_n22879), .O(new_n22932));
  nor2 g22739(.a(new_n22873), .b(new_n22867), .O(new_n22933));
  inv1 g22740(.a(new_n22933), .O(new_n22934));
  nor2 g22741(.a(new_n10895), .b(new_n8476), .O(new_n22935));
  inv1 g22742(.a(new_n22935), .O(new_n22936));
  nor2 g22743(.a(new_n10468), .b(new_n8946), .O(new_n22937));
  nor2 g22744(.a(new_n22937), .b(new_n22900), .O(new_n22938));
  nor2 g22745(.a(new_n10468), .b(new_n9156), .O(new_n22939));
  inv1 g22746(.a(new_n22939), .O(new_n22940));
  nor2 g22747(.a(new_n22940), .b(new_n22814), .O(new_n22941));
  nor2 g22748(.a(new_n22941), .b(new_n22938), .O(new_n22942));
  nor2 g22749(.a(new_n22942), .b(new_n22936), .O(new_n22943));
  inv1 g22750(.a(new_n22942), .O(new_n22944));
  nor2 g22751(.a(new_n22944), .b(new_n22935), .O(new_n22945));
  nor2 g22752(.a(new_n22945), .b(new_n22943), .O(new_n22946));
  nor2 g22753(.a(new_n9873), .b(\a[57] ), .O(new_n22947));
  nor2 g22754(.a(new_n22947), .b(new_n22888), .O(new_n22948));
  inv1 g22755(.a(new_n22947), .O(new_n22949));
  nor2 g22756(.a(new_n22949), .b(new_n22887), .O(new_n22950));
  nor2 g22757(.a(new_n22950), .b(new_n22948), .O(new_n22951));
  nor2 g22758(.a(new_n22951), .b(new_n22946), .O(new_n22952));
  inv1 g22759(.a(new_n22946), .O(new_n22953));
  inv1 g22760(.a(new_n22951), .O(new_n22954));
  nor2 g22761(.a(new_n22954), .b(new_n22953), .O(new_n22955));
  nor2 g22762(.a(new_n22955), .b(new_n22952), .O(new_n22956));
  nor2 g22763(.a(new_n22956), .b(new_n22934), .O(new_n22957));
  inv1 g22764(.a(new_n22956), .O(new_n22958));
  nor2 g22765(.a(new_n22958), .b(new_n22933), .O(new_n22959));
  nor2 g22766(.a(new_n22959), .b(new_n22957), .O(new_n22960));
  inv1 g22767(.a(new_n22960), .O(new_n22961));
  nor2 g22768(.a(new_n11596), .b(new_n8026), .O(new_n22962));
  inv1 g22769(.a(new_n22962), .O(new_n22963));
  nor2 g22770(.a(new_n22906), .b(new_n22899), .O(new_n22964));
  inv1 g22771(.a(new_n22964), .O(new_n22965));
  nor2 g22772(.a(new_n22965), .b(new_n22963), .O(new_n22966));
  nor2 g22773(.a(new_n22964), .b(new_n22962), .O(new_n22967));
  nor2 g22774(.a(new_n22967), .b(new_n22966), .O(new_n22968));
  nor2 g22775(.a(new_n22892), .b(new_n22886), .O(new_n22969));
  nor2 g22776(.a(new_n22969), .b(new_n22968), .O(new_n22970));
  inv1 g22777(.a(new_n22968), .O(new_n22971));
  inv1 g22778(.a(new_n22969), .O(new_n22972));
  nor2 g22779(.a(new_n22972), .b(new_n22971), .O(new_n22973));
  nor2 g22780(.a(new_n22973), .b(new_n22970), .O(new_n22974));
  nor2 g22781(.a(new_n22915), .b(new_n22908), .O(new_n22975));
  inv1 g22782(.a(new_n22975), .O(new_n22976));
  nor2 g22783(.a(new_n22976), .b(new_n22974), .O(new_n22977));
  inv1 g22784(.a(new_n22974), .O(new_n22978));
  nor2 g22785(.a(new_n22975), .b(new_n22978), .O(new_n22979));
  nor2 g22786(.a(new_n22979), .b(new_n22977), .O(new_n22980));
  inv1 g22787(.a(new_n22980), .O(new_n22981));
  nor2 g22788(.a(new_n22981), .b(new_n22961), .O(new_n22982));
  nor2 g22789(.a(new_n22980), .b(new_n22960), .O(new_n22983));
  nor2 g22790(.a(new_n22983), .b(new_n22982), .O(new_n22984));
  inv1 g22791(.a(new_n22984), .O(new_n22985));
  nor2 g22792(.a(new_n22985), .b(new_n22932), .O(new_n22986));
  inv1 g22793(.a(new_n22932), .O(new_n22987));
  nor2 g22794(.a(new_n22984), .b(new_n22987), .O(new_n22988));
  nor2 g22795(.a(new_n22988), .b(new_n22986), .O(new_n22989));
  inv1 g22796(.a(new_n22989), .O(new_n22990));
  nor2 g22797(.a(new_n22928), .b(new_n22923), .O(new_n22991));
  inv1 g22798(.a(new_n22991), .O(new_n22992));
  nor2 g22799(.a(new_n22992), .b(new_n22990), .O(new_n22993));
  nor2 g22800(.a(new_n22991), .b(new_n22989), .O(new_n22994));
  nor2 g22801(.a(new_n22994), .b(new_n22993), .O(new_n22995));
  inv1 g22802(.a(new_n22995), .O(\asquared[116] ));
  nor2 g22803(.a(new_n22959), .b(new_n22952), .O(new_n22997));
  inv1 g22804(.a(new_n22997), .O(new_n22998));
  nor2 g22805(.a(new_n22973), .b(new_n22966), .O(new_n22999));
  inv1 g22806(.a(new_n22999), .O(new_n23000));
  nor2 g22807(.a(new_n23000), .b(new_n22998), .O(new_n23001));
  nor2 g22808(.a(new_n22999), .b(new_n22997), .O(new_n23002));
  nor2 g22809(.a(new_n23002), .b(new_n23001), .O(new_n23003));
  inv1 g22810(.a(new_n23003), .O(new_n23004));
  nor2 g22811(.a(new_n11186), .b(new_n8476), .O(new_n23005));
  nor2 g22812(.a(new_n11596), .b(new_n8170), .O(new_n23006));
  nor2 g22813(.a(new_n23006), .b(new_n23005), .O(new_n23007));
  nor2 g22814(.a(new_n11596), .b(new_n8476), .O(new_n23008));
  inv1 g22815(.a(new_n23008), .O(new_n23009));
  nor2 g22816(.a(new_n23009), .b(new_n22888), .O(new_n23010));
  nor2 g22817(.a(new_n23010), .b(new_n23007), .O(new_n23011));
  inv1 g22818(.a(new_n23011), .O(new_n23012));
  nor2 g22819(.a(new_n22950), .b(new_n9873), .O(new_n23013));
  inv1 g22820(.a(new_n23013), .O(new_n23014));
  nor2 g22821(.a(new_n23014), .b(new_n23012), .O(new_n23015));
  nor2 g22822(.a(new_n23013), .b(new_n23011), .O(new_n23016));
  nor2 g22823(.a(new_n23016), .b(new_n23015), .O(new_n23017));
  inv1 g22824(.a(new_n23017), .O(new_n23018));
  nor2 g22825(.a(new_n10895), .b(new_n8946), .O(new_n23019));
  inv1 g22826(.a(new_n23019), .O(new_n23020));
  nor2 g22827(.a(new_n10320), .b(new_n9658), .O(new_n23021));
  nor2 g22828(.a(new_n23021), .b(new_n22939), .O(new_n23022));
  nor2 g22829(.a(new_n10468), .b(new_n9658), .O(new_n23023));
  inv1 g22830(.a(new_n23023), .O(new_n23024));
  nor2 g22831(.a(new_n23024), .b(new_n22901), .O(new_n23025));
  nor2 g22832(.a(new_n23025), .b(new_n23022), .O(new_n23026));
  nor2 g22833(.a(new_n23026), .b(new_n23020), .O(new_n23027));
  inv1 g22834(.a(new_n23026), .O(new_n23028));
  nor2 g22835(.a(new_n23028), .b(new_n23019), .O(new_n23029));
  nor2 g22836(.a(new_n23029), .b(new_n23027), .O(new_n23030));
  nor2 g22837(.a(new_n22945), .b(new_n22938), .O(new_n23031));
  inv1 g22838(.a(new_n23031), .O(new_n23032));
  nor2 g22839(.a(new_n23032), .b(new_n23030), .O(new_n23033));
  inv1 g22840(.a(new_n23030), .O(new_n23034));
  nor2 g22841(.a(new_n23031), .b(new_n23034), .O(new_n23035));
  nor2 g22842(.a(new_n23035), .b(new_n23033), .O(new_n23036));
  inv1 g22843(.a(new_n23036), .O(new_n23037));
  nor2 g22844(.a(new_n23037), .b(new_n23018), .O(new_n23038));
  nor2 g22845(.a(new_n23036), .b(new_n23017), .O(new_n23039));
  nor2 g22846(.a(new_n23039), .b(new_n23038), .O(new_n23040));
  inv1 g22847(.a(new_n23040), .O(new_n23041));
  nor2 g22848(.a(new_n23041), .b(new_n23004), .O(new_n23042));
  nor2 g22849(.a(new_n23040), .b(new_n23003), .O(new_n23043));
  nor2 g22850(.a(new_n23043), .b(new_n23042), .O(new_n23044));
  nor2 g22851(.a(new_n22982), .b(new_n22979), .O(new_n23045));
  inv1 g22852(.a(new_n23045), .O(new_n23046));
  nor2 g22853(.a(new_n23046), .b(new_n23044), .O(new_n23047));
  inv1 g22854(.a(new_n23044), .O(new_n23048));
  nor2 g22855(.a(new_n23045), .b(new_n23048), .O(new_n23049));
  nor2 g22856(.a(new_n23049), .b(new_n23047), .O(new_n23050));
  inv1 g22857(.a(new_n23050), .O(new_n23051));
  nor2 g22858(.a(new_n22991), .b(new_n22988), .O(new_n23052));
  nor2 g22859(.a(new_n23052), .b(new_n22986), .O(new_n23053));
  nor2 g22860(.a(new_n23053), .b(new_n23051), .O(new_n23054));
  inv1 g22861(.a(new_n23053), .O(new_n23055));
  nor2 g22862(.a(new_n23055), .b(new_n23050), .O(new_n23056));
  nor2 g22863(.a(new_n23056), .b(new_n23054), .O(\asquared[117] ));
  nor2 g22864(.a(new_n23042), .b(new_n23002), .O(new_n23058));
  nor2 g22865(.a(new_n23038), .b(new_n23033), .O(new_n23059));
  nor2 g22866(.a(new_n11186), .b(new_n8946), .O(new_n23060));
  inv1 g22867(.a(new_n23060), .O(new_n23061));
  nor2 g22868(.a(new_n10320), .b(\a[58] ), .O(new_n23062));
  nor2 g22869(.a(new_n23062), .b(new_n23061), .O(new_n23063));
  inv1 g22870(.a(new_n23062), .O(new_n23064));
  nor2 g22871(.a(new_n23064), .b(new_n23060), .O(new_n23065));
  nor2 g22872(.a(new_n23065), .b(new_n23063), .O(new_n23066));
  nor2 g22873(.a(new_n23066), .b(new_n23059), .O(new_n23067));
  inv1 g22874(.a(new_n23059), .O(new_n23068));
  inv1 g22875(.a(new_n23066), .O(new_n23069));
  nor2 g22876(.a(new_n23069), .b(new_n23068), .O(new_n23070));
  nor2 g22877(.a(new_n23070), .b(new_n23067), .O(new_n23071));
  inv1 g22878(.a(new_n23071), .O(new_n23072));
  nor2 g22879(.a(new_n23015), .b(new_n23010), .O(new_n23073));
  inv1 g22880(.a(new_n23073), .O(new_n23074));
  nor2 g22881(.a(new_n23029), .b(new_n23022), .O(new_n23075));
  nor2 g22882(.a(new_n23075), .b(new_n23074), .O(new_n23076));
  inv1 g22883(.a(new_n23075), .O(new_n23077));
  nor2 g22884(.a(new_n23077), .b(new_n23073), .O(new_n23078));
  nor2 g22885(.a(new_n23078), .b(new_n23076), .O(new_n23079));
  inv1 g22886(.a(new_n23079), .O(new_n23080));
  nor2 g22887(.a(new_n10895), .b(new_n9156), .O(new_n23081));
  nor2 g22888(.a(new_n23081), .b(new_n23023), .O(new_n23082));
  nor2 g22889(.a(new_n10895), .b(new_n9658), .O(new_n23083));
  inv1 g22890(.a(new_n23083), .O(new_n23084));
  nor2 g22891(.a(new_n23084), .b(new_n22940), .O(new_n23085));
  nor2 g22892(.a(new_n23085), .b(new_n23082), .O(new_n23086));
  nor2 g22893(.a(new_n23086), .b(new_n23009), .O(new_n23087));
  inv1 g22894(.a(new_n23086), .O(new_n23088));
  nor2 g22895(.a(new_n23088), .b(new_n23008), .O(new_n23089));
  nor2 g22896(.a(new_n23089), .b(new_n23087), .O(new_n23090));
  nor2 g22897(.a(new_n23090), .b(new_n23080), .O(new_n23091));
  inv1 g22898(.a(new_n23090), .O(new_n23092));
  nor2 g22899(.a(new_n23092), .b(new_n23079), .O(new_n23093));
  nor2 g22900(.a(new_n23093), .b(new_n23091), .O(new_n23094));
  inv1 g22901(.a(new_n23094), .O(new_n23095));
  nor2 g22902(.a(new_n23095), .b(new_n23072), .O(new_n23096));
  nor2 g22903(.a(new_n23094), .b(new_n23071), .O(new_n23097));
  nor2 g22904(.a(new_n23097), .b(new_n23096), .O(new_n23098));
  inv1 g22905(.a(new_n23098), .O(new_n23099));
  nor2 g22906(.a(new_n23099), .b(new_n23058), .O(new_n23100));
  inv1 g22907(.a(new_n23058), .O(new_n23101));
  nor2 g22908(.a(new_n23098), .b(new_n23101), .O(new_n23102));
  nor2 g22909(.a(new_n23102), .b(new_n23100), .O(new_n23103));
  inv1 g22910(.a(new_n23103), .O(new_n23104));
  nor2 g22911(.a(new_n23054), .b(new_n23049), .O(new_n23105));
  inv1 g22912(.a(new_n23105), .O(new_n23106));
  nor2 g22913(.a(new_n23106), .b(new_n23104), .O(new_n23107));
  nor2 g22914(.a(new_n23105), .b(new_n23103), .O(new_n23108));
  nor2 g22915(.a(new_n23108), .b(new_n23107), .O(new_n23109));
  inv1 g22916(.a(new_n23109), .O(\asquared[118] ));
  nor2 g22917(.a(new_n11596), .b(new_n8946), .O(new_n23111));
  inv1 g22918(.a(new_n23111), .O(new_n23112));
  nor2 g22919(.a(new_n23065), .b(new_n10320), .O(new_n23113));
  inv1 g22920(.a(new_n23113), .O(new_n23114));
  nor2 g22921(.a(new_n23114), .b(new_n23112), .O(new_n23115));
  nor2 g22922(.a(new_n23113), .b(new_n23111), .O(new_n23116));
  nor2 g22923(.a(new_n23116), .b(new_n23115), .O(new_n23117));
  nor2 g22924(.a(new_n23089), .b(new_n23082), .O(new_n23118));
  nor2 g22925(.a(new_n23118), .b(new_n23117), .O(new_n23119));
  inv1 g22926(.a(new_n23117), .O(new_n23120));
  inv1 g22927(.a(new_n23118), .O(new_n23121));
  nor2 g22928(.a(new_n23121), .b(new_n23120), .O(new_n23122));
  nor2 g22929(.a(new_n23122), .b(new_n23119), .O(new_n23123));
  nor2 g22930(.a(new_n11186), .b(new_n9156), .O(new_n23124));
  inv1 g22931(.a(new_n23124), .O(new_n23125));
  nor2 g22932(.a(new_n10468), .b(new_n9873), .O(new_n23126));
  nor2 g22933(.a(new_n23126), .b(new_n23083), .O(new_n23127));
  nor2 g22934(.a(new_n10895), .b(new_n9873), .O(new_n23128));
  inv1 g22935(.a(new_n23128), .O(new_n23129));
  nor2 g22936(.a(new_n23129), .b(new_n23024), .O(new_n23130));
  nor2 g22937(.a(new_n23130), .b(new_n23127), .O(new_n23131));
  nor2 g22938(.a(new_n23131), .b(new_n23125), .O(new_n23132));
  inv1 g22939(.a(new_n23131), .O(new_n23133));
  nor2 g22940(.a(new_n23133), .b(new_n23124), .O(new_n23134));
  nor2 g22941(.a(new_n23134), .b(new_n23132), .O(new_n23135));
  nor2 g22942(.a(new_n23091), .b(new_n23078), .O(new_n23136));
  nor2 g22943(.a(new_n23136), .b(new_n23135), .O(new_n23137));
  inv1 g22944(.a(new_n23135), .O(new_n23138));
  inv1 g22945(.a(new_n23136), .O(new_n23139));
  nor2 g22946(.a(new_n23139), .b(new_n23138), .O(new_n23140));
  nor2 g22947(.a(new_n23140), .b(new_n23137), .O(new_n23141));
  nor2 g22948(.a(new_n23141), .b(new_n23123), .O(new_n23142));
  inv1 g22949(.a(new_n23123), .O(new_n23143));
  inv1 g22950(.a(new_n23141), .O(new_n23144));
  nor2 g22951(.a(new_n23144), .b(new_n23143), .O(new_n23145));
  nor2 g22952(.a(new_n23145), .b(new_n23142), .O(new_n23146));
  nor2 g22953(.a(new_n23096), .b(new_n23067), .O(new_n23147));
  inv1 g22954(.a(new_n23147), .O(new_n23148));
  nor2 g22955(.a(new_n23148), .b(new_n23146), .O(new_n23149));
  inv1 g22956(.a(new_n23146), .O(new_n23150));
  nor2 g22957(.a(new_n23147), .b(new_n23150), .O(new_n23151));
  nor2 g22958(.a(new_n23151), .b(new_n23149), .O(new_n23152));
  inv1 g22959(.a(new_n23152), .O(new_n23153));
  nor2 g22960(.a(new_n23105), .b(new_n23102), .O(new_n23154));
  nor2 g22961(.a(new_n23154), .b(new_n23100), .O(new_n23155));
  nor2 g22962(.a(new_n23155), .b(new_n23153), .O(new_n23156));
  inv1 g22963(.a(new_n23155), .O(new_n23157));
  nor2 g22964(.a(new_n23157), .b(new_n23152), .O(new_n23158));
  nor2 g22965(.a(new_n23158), .b(new_n23156), .O(\asquared[119] ));
  nor2 g22966(.a(new_n23122), .b(new_n23115), .O(new_n23160));
  inv1 g22967(.a(new_n23160), .O(new_n23161));
  nor2 g22968(.a(new_n11596), .b(new_n9156), .O(new_n23162));
  nor2 g22969(.a(new_n23162), .b(new_n23128), .O(new_n23163));
  inv1 g22970(.a(new_n23081), .O(new_n23164));
  nor2 g22971(.a(new_n11596), .b(new_n9873), .O(new_n23165));
  inv1 g22972(.a(new_n23165), .O(new_n23166));
  nor2 g22973(.a(new_n23166), .b(new_n23164), .O(new_n23167));
  nor2 g22974(.a(new_n23167), .b(new_n23163), .O(new_n23168));
  inv1 g22975(.a(new_n23168), .O(new_n23169));
  nor2 g22976(.a(new_n23134), .b(new_n23127), .O(new_n23170));
  inv1 g22977(.a(new_n23170), .O(new_n23171));
  nor2 g22978(.a(new_n23171), .b(new_n23169), .O(new_n23172));
  nor2 g22979(.a(new_n23170), .b(new_n23168), .O(new_n23173));
  nor2 g22980(.a(new_n23173), .b(new_n23172), .O(new_n23174));
  inv1 g22981(.a(new_n23174), .O(new_n23175));
  nor2 g22982(.a(new_n11186), .b(new_n9658), .O(new_n23176));
  inv1 g22983(.a(new_n23176), .O(new_n23177));
  nor2 g22984(.a(new_n10468), .b(\a[59] ), .O(new_n23178));
  nor2 g22985(.a(new_n23178), .b(new_n23177), .O(new_n23179));
  inv1 g22986(.a(new_n23178), .O(new_n23180));
  nor2 g22987(.a(new_n23180), .b(new_n23176), .O(new_n23181));
  nor2 g22988(.a(new_n23181), .b(new_n23179), .O(new_n23182));
  nor2 g22989(.a(new_n23182), .b(new_n23175), .O(new_n23183));
  inv1 g22990(.a(new_n23182), .O(new_n23184));
  nor2 g22991(.a(new_n23184), .b(new_n23174), .O(new_n23185));
  nor2 g22992(.a(new_n23185), .b(new_n23183), .O(new_n23186));
  nor2 g22993(.a(new_n23186), .b(new_n23161), .O(new_n23187));
  inv1 g22994(.a(new_n23186), .O(new_n23188));
  nor2 g22995(.a(new_n23188), .b(new_n23160), .O(new_n23189));
  nor2 g22996(.a(new_n23189), .b(new_n23187), .O(new_n23190));
  inv1 g22997(.a(new_n23190), .O(new_n23191));
  nor2 g22998(.a(new_n23145), .b(new_n23137), .O(new_n23192));
  nor2 g22999(.a(new_n23192), .b(new_n23191), .O(new_n23193));
  inv1 g23000(.a(new_n23192), .O(new_n23194));
  nor2 g23001(.a(new_n23194), .b(new_n23190), .O(new_n23195));
  nor2 g23002(.a(new_n23195), .b(new_n23193), .O(new_n23196));
  inv1 g23003(.a(new_n23196), .O(new_n23197));
  nor2 g23004(.a(new_n23156), .b(new_n23151), .O(new_n23198));
  nor2 g23005(.a(new_n23198), .b(new_n23197), .O(new_n23199));
  inv1 g23006(.a(new_n23198), .O(new_n23200));
  nor2 g23007(.a(new_n23200), .b(new_n23196), .O(new_n23201));
  nor2 g23008(.a(new_n23201), .b(new_n23199), .O(\asquared[120] ));
  nor2 g23009(.a(new_n23189), .b(new_n23183), .O(new_n23203));
  inv1 g23010(.a(new_n23203), .O(new_n23204));
  nor2 g23011(.a(new_n23172), .b(new_n23167), .O(new_n23205));
  inv1 g23012(.a(new_n23205), .O(new_n23206));
  nor2 g23013(.a(new_n23181), .b(new_n10468), .O(new_n23207));
  nor2 g23014(.a(new_n23207), .b(new_n23206), .O(new_n23208));
  inv1 g23015(.a(new_n23207), .O(new_n23209));
  nor2 g23016(.a(new_n23209), .b(new_n23205), .O(new_n23210));
  nor2 g23017(.a(new_n23210), .b(new_n23208), .O(new_n23211));
  inv1 g23018(.a(new_n23211), .O(new_n23212));
  nor2 g23019(.a(new_n11596), .b(new_n9658), .O(new_n23213));
  inv1 g23020(.a(new_n23213), .O(new_n23214));
  nor2 g23021(.a(new_n11186), .b(new_n9873), .O(new_n23215));
  nor2 g23022(.a(new_n10895), .b(new_n10320), .O(new_n23216));
  nor2 g23023(.a(new_n23216), .b(new_n23215), .O(new_n23217));
  nor2 g23024(.a(new_n11186), .b(new_n10320), .O(new_n23218));
  inv1 g23025(.a(new_n23218), .O(new_n23219));
  nor2 g23026(.a(new_n23219), .b(new_n23129), .O(new_n23220));
  nor2 g23027(.a(new_n23220), .b(new_n23217), .O(new_n23221));
  nor2 g23028(.a(new_n23221), .b(new_n23214), .O(new_n23222));
  inv1 g23029(.a(new_n23221), .O(new_n23223));
  nor2 g23030(.a(new_n23223), .b(new_n23213), .O(new_n23224));
  nor2 g23031(.a(new_n23224), .b(new_n23222), .O(new_n23225));
  nor2 g23032(.a(new_n23225), .b(new_n23212), .O(new_n23226));
  inv1 g23033(.a(new_n23225), .O(new_n23227));
  nor2 g23034(.a(new_n23227), .b(new_n23211), .O(new_n23228));
  nor2 g23035(.a(new_n23228), .b(new_n23226), .O(new_n23229));
  nor2 g23036(.a(new_n23229), .b(new_n23204), .O(new_n23230));
  inv1 g23037(.a(new_n23229), .O(new_n23231));
  nor2 g23038(.a(new_n23231), .b(new_n23203), .O(new_n23232));
  nor2 g23039(.a(new_n23232), .b(new_n23230), .O(new_n23233));
  inv1 g23040(.a(new_n23233), .O(new_n23234));
  nor2 g23041(.a(new_n23199), .b(new_n23193), .O(new_n23235));
  nor2 g23042(.a(new_n23235), .b(new_n23234), .O(new_n23236));
  inv1 g23043(.a(new_n23235), .O(new_n23237));
  nor2 g23044(.a(new_n23237), .b(new_n23233), .O(new_n23238));
  nor2 g23045(.a(new_n23238), .b(new_n23236), .O(\asquared[121] ));
  nor2 g23046(.a(new_n23224), .b(new_n23217), .O(new_n23240));
  inv1 g23047(.a(new_n23240), .O(new_n23241));
  nor2 g23048(.a(new_n23241), .b(new_n23166), .O(new_n23242));
  nor2 g23049(.a(new_n23240), .b(new_n23165), .O(new_n23243));
  nor2 g23050(.a(new_n23243), .b(new_n23242), .O(new_n23244));
  nor2 g23051(.a(new_n10895), .b(\a[60] ), .O(new_n23245));
  nor2 g23052(.a(new_n23245), .b(new_n23219), .O(new_n23246));
  inv1 g23053(.a(new_n23245), .O(new_n23247));
  nor2 g23054(.a(new_n23247), .b(new_n23218), .O(new_n23248));
  nor2 g23055(.a(new_n23248), .b(new_n23246), .O(new_n23249));
  inv1 g23056(.a(new_n23249), .O(new_n23250));
  nor2 g23057(.a(new_n23250), .b(new_n23244), .O(new_n23251));
  inv1 g23058(.a(new_n23244), .O(new_n23252));
  nor2 g23059(.a(new_n23249), .b(new_n23252), .O(new_n23253));
  nor2 g23060(.a(new_n23253), .b(new_n23251), .O(new_n23254));
  nor2 g23061(.a(new_n23226), .b(new_n23210), .O(new_n23255));
  inv1 g23062(.a(new_n23255), .O(new_n23256));
  nor2 g23063(.a(new_n23256), .b(new_n23254), .O(new_n23257));
  inv1 g23064(.a(new_n23254), .O(new_n23258));
  nor2 g23065(.a(new_n23255), .b(new_n23258), .O(new_n23259));
  nor2 g23066(.a(new_n23259), .b(new_n23257), .O(new_n23260));
  inv1 g23067(.a(new_n23260), .O(new_n23261));
  nor2 g23068(.a(new_n23236), .b(new_n23232), .O(new_n23262));
  nor2 g23069(.a(new_n23262), .b(new_n23261), .O(new_n23263));
  inv1 g23070(.a(new_n23262), .O(new_n23264));
  nor2 g23071(.a(new_n23264), .b(new_n23260), .O(new_n23265));
  nor2 g23072(.a(new_n23265), .b(new_n23263), .O(\asquared[122] ));
  nor2 g23073(.a(new_n23253), .b(new_n23242), .O(new_n23267));
  inv1 g23074(.a(new_n23267), .O(new_n23268));
  nor2 g23075(.a(new_n11186), .b(new_n10468), .O(new_n23269));
  nor2 g23076(.a(new_n11596), .b(new_n10320), .O(new_n23270));
  nor2 g23077(.a(new_n23270), .b(new_n23269), .O(new_n23271));
  nor2 g23078(.a(new_n11596), .b(new_n10468), .O(new_n23272));
  inv1 g23079(.a(new_n23272), .O(new_n23273));
  nor2 g23080(.a(new_n23273), .b(new_n23219), .O(new_n23274));
  nor2 g23081(.a(new_n23274), .b(new_n23271), .O(new_n23275));
  inv1 g23082(.a(new_n23275), .O(new_n23276));
  nor2 g23083(.a(new_n23248), .b(new_n10895), .O(new_n23277));
  inv1 g23084(.a(new_n23277), .O(new_n23278));
  nor2 g23085(.a(new_n23278), .b(new_n23276), .O(new_n23279));
  nor2 g23086(.a(new_n23277), .b(new_n23275), .O(new_n23280));
  nor2 g23087(.a(new_n23280), .b(new_n23279), .O(new_n23281));
  nor2 g23088(.a(new_n23281), .b(new_n23268), .O(new_n23282));
  inv1 g23089(.a(new_n23281), .O(new_n23283));
  nor2 g23090(.a(new_n23283), .b(new_n23267), .O(new_n23284));
  nor2 g23091(.a(new_n23284), .b(new_n23282), .O(new_n23285));
  inv1 g23092(.a(new_n23285), .O(new_n23286));
  nor2 g23093(.a(new_n23263), .b(new_n23259), .O(new_n23287));
  nor2 g23094(.a(new_n23287), .b(new_n23286), .O(new_n23288));
  inv1 g23095(.a(new_n23287), .O(new_n23289));
  nor2 g23096(.a(new_n23289), .b(new_n23285), .O(new_n23290));
  nor2 g23097(.a(new_n23290), .b(new_n23288), .O(\asquared[123] ));
  nor2 g23098(.a(new_n23279), .b(new_n23274), .O(new_n23292));
  inv1 g23099(.a(new_n23292), .O(new_n23293));
  nor2 g23100(.a(new_n11186), .b(\a[61] ), .O(new_n23294));
  inv1 g23101(.a(new_n23294), .O(new_n23295));
  nor2 g23102(.a(new_n23295), .b(new_n23272), .O(new_n23296));
  nor2 g23103(.a(new_n23294), .b(new_n23273), .O(new_n23297));
  nor2 g23104(.a(new_n23297), .b(new_n23296), .O(new_n23298));
  inv1 g23105(.a(new_n23298), .O(new_n23299));
  nor2 g23106(.a(new_n23299), .b(new_n23293), .O(new_n23300));
  nor2 g23107(.a(new_n23298), .b(new_n23292), .O(new_n23301));
  nor2 g23108(.a(new_n23301), .b(new_n23300), .O(new_n23302));
  inv1 g23109(.a(new_n23302), .O(new_n23303));
  nor2 g23110(.a(new_n23288), .b(new_n23284), .O(new_n23304));
  nor2 g23111(.a(new_n23304), .b(new_n23303), .O(new_n23305));
  inv1 g23112(.a(new_n23304), .O(new_n23306));
  nor2 g23113(.a(new_n23306), .b(new_n23302), .O(new_n23307));
  nor2 g23114(.a(new_n23307), .b(new_n23305), .O(\asquared[124] ));
  nor2 g23115(.a(new_n11596), .b(new_n10895), .O(new_n23309));
  inv1 g23116(.a(new_n23309), .O(new_n23310));
  nor2 g23117(.a(new_n23310), .b(new_n11186), .O(new_n23311));
  nor2 g23118(.a(new_n23299), .b(new_n11186), .O(new_n23312));
  nor2 g23119(.a(new_n23312), .b(new_n23309), .O(new_n23313));
  nor2 g23120(.a(new_n23313), .b(new_n23311), .O(new_n23314));
  nor2 g23121(.a(new_n23305), .b(new_n23301), .O(new_n23315));
  inv1 g23122(.a(new_n23315), .O(new_n23316));
  nor2 g23123(.a(new_n23316), .b(new_n23314), .O(new_n23317));
  inv1 g23124(.a(new_n23314), .O(new_n23318));
  nor2 g23125(.a(new_n23315), .b(new_n23318), .O(new_n23319));
  nor2 g23126(.a(new_n23319), .b(new_n23317), .O(\asquared[125] ));
  nor2 g23127(.a(new_n23315), .b(new_n23313), .O(new_n23321));
  nor2 g23128(.a(new_n23294), .b(new_n11596), .O(new_n23322));
  nor2 g23129(.a(new_n23322), .b(new_n23321), .O(new_n23323));
  inv1 g23130(.a(new_n23321), .O(new_n23324));
  nor2 g23131(.a(new_n11596), .b(\a[62] ), .O(new_n23325));
  inv1 g23132(.a(new_n23325), .O(new_n23326));
  nor2 g23133(.a(new_n23326), .b(new_n23324), .O(new_n23327));
  nor2 g23134(.a(new_n23327), .b(new_n23323), .O(\asquared[126] ));
  nor2 g23135(.a(new_n23321), .b(\a[62] ), .O(new_n23329));
  nor2 g23136(.a(new_n23329), .b(new_n11596), .O(\asquared[127] ));
  zero g23137(.O(\asquared[1] ));
  buf  g23138(.a(\a[0] ), .O(\asquared[0] ));
endmodule


