// Benchmark "top" written by ABC on Tue Nov 26 20:40:42 2024

module top ( 
    _9, _8, _7, _6, _5, _4, _3, _2, _1,
    _52  );
  input  _9, _8, _7, _6, _5, _4, _3, _2, _1;
  output _52;
  wire new_n11, new_n12, new_n13, new_n14, new_n15, new_n16, new_n17,
    new_n18, new_n19, new_n20, new_n21, new_n22, new_n23, new_n24, new_n25,
    new_n26, new_n27, new_n28, new_n29, new_n30, new_n31, new_n32, new_n33,
    new_n34, new_n35, new_n36, new_n37, new_n38, new_n39, new_n40, new_n41,
    new_n42, new_n43, new_n44, new_n45, new_n46, new_n47, new_n48, new_n49,
    new_n50, new_n51, new_n52, new_n53, new_n54, new_n55, new_n56, new_n57,
    new_n58, new_n59, new_n60, new_n61, new_n62, new_n63, new_n64, new_n65,
    new_n66, new_n67, new_n68, new_n69, new_n70, new_n71, new_n72, new_n73,
    new_n74, new_n75, new_n76, new_n77, new_n78, new_n79, new_n80, new_n81,
    new_n82, new_n83, new_n84, new_n85, new_n86, new_n87, new_n88, new_n89,
    new_n90, new_n91, new_n92, new_n93, new_n94, new_n95, new_n96, new_n97,
    new_n98, new_n99, new_n100, new_n101, new_n102, new_n103, new_n104,
    new_n105, new_n106, new_n107, new_n108, new_n109, new_n110, new_n111,
    new_n112, new_n113, new_n114, new_n115, new_n116, new_n117, new_n118,
    new_n119, new_n120, new_n121, new_n122, new_n123, new_n124, new_n125,
    new_n126, new_n127, new_n128, new_n129, new_n130, new_n131, new_n132,
    new_n133, new_n134, new_n135, new_n136, new_n137, new_n138, new_n139,
    new_n140, new_n141, new_n142, new_n143, new_n144, new_n145, new_n146,
    new_n147, new_n148, new_n149, new_n150, new_n151, new_n152, new_n153,
    new_n154, new_n155, new_n156, new_n157, new_n158, new_n159, new_n160,
    new_n161, new_n162, new_n163, new_n164, new_n165, new_n166, new_n167,
    new_n168, new_n169, new_n170, new_n171, new_n172, new_n173, new_n174,
    new_n175, new_n176, new_n177, new_n178, new_n179, new_n180, new_n181,
    new_n182, new_n183, new_n184, new_n185, new_n186, new_n187, new_n188,
    new_n189, new_n190, new_n191, new_n192, new_n193, new_n194, new_n195,
    new_n196, new_n197, new_n198, new_n199, new_n200, new_n201, new_n202,
    new_n203, new_n204, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n235, new_n236, new_n237,
    new_n238, new_n239, new_n240, new_n241, new_n242, new_n243, new_n244,
    new_n245, new_n246, new_n247, new_n248, new_n249, new_n250, new_n251,
    new_n252, new_n253, new_n254, new_n255, new_n256, new_n257, new_n258,
    new_n259, new_n260, new_n261, new_n262, new_n263, new_n264, new_n265,
    new_n266, new_n267, new_n268, new_n269, new_n270, new_n271, new_n272,
    new_n273, new_n274, new_n275, new_n276, new_n277, new_n278, new_n279;
  inv1 g000(.a(_8), .O(new_n11));
  inv1 g001(.a(_7), .O(new_n12));
  inv1 g002(.a(_6), .O(new_n13));
  nor2 g003(.a(_2), .b(new_n13), .O(new_n14));
  inv1 g004(.a(_3), .O(new_n15));
  nor2 g005(.a(new_n15), .b(_4), .O(new_n16));
  nor2 g006(.a(new_n16), .b(new_n14), .O(new_n17));
  nor2 g007(.a(new_n17), .b(new_n12), .O(new_n18));
  inv1 g008(.a(_5), .O(new_n19));
  inv1 g009(.a(_4), .O(new_n20));
  nor2 g010(.a(_3), .b(new_n20), .O(new_n21));
  inv1 g011(.a(new_n21), .O(new_n22));
  nor2 g012(.a(new_n22), .b(new_n19), .O(new_n23));
  nor2 g013(.a(new_n15), .b(_5), .O(new_n24));
  nor2 g014(.a(new_n20), .b(_7), .O(new_n25));
  nor2 g015(.a(new_n25), .b(new_n24), .O(new_n26));
  nor2 g016(.a(new_n26), .b(new_n13), .O(new_n27));
  nor2 g017(.a(new_n27), .b(new_n23), .O(new_n28));
  inv1 g018(.a(new_n28), .O(new_n29));
  nor2 g019(.a(new_n29), .b(new_n18), .O(new_n30));
  nor2 g020(.a(new_n30), .b(_9), .O(new_n31));
  inv1 g021(.a(_9), .O(new_n32));
  nor2 g022(.a(_3), .b(new_n32), .O(new_n33));
  inv1 g023(.a(new_n33), .O(new_n34));
  nor2 g024(.a(_2), .b(new_n12), .O(new_n35));
  inv1 g025(.a(new_n35), .O(new_n36));
  nor2 g026(.a(new_n36), .b(new_n34), .O(new_n37));
  nor2 g027(.a(new_n19), .b(_7), .O(new_n38));
  nor2 g028(.a(_5), .b(new_n32), .O(new_n39));
  nor2 g029(.a(new_n39), .b(new_n38), .O(new_n40));
  nor2 g030(.a(new_n15), .b(_6), .O(new_n41));
  inv1 g031(.a(new_n41), .O(new_n42));
  nor2 g032(.a(new_n42), .b(new_n40), .O(new_n43));
  nor2 g033(.a(new_n43), .b(new_n37), .O(new_n44));
  inv1 g034(.a(new_n44), .O(new_n45));
  nor2 g035(.a(new_n45), .b(new_n31), .O(new_n46));
  nor2 g036(.a(new_n46), .b(new_n11), .O(new_n47));
  inv1 g037(.a(new_n24), .O(new_n48));
  inv1 g038(.a(_2), .O(new_n49));
  inv1 g039(.a(new_n25), .O(new_n50));
  nor2 g040(.a(new_n50), .b(new_n49), .O(new_n51));
  nor2 g041(.a(_8), .b(new_n32), .O(new_n52));
  inv1 g042(.a(new_n52), .O(new_n53));
  nor2 g043(.a(new_n53), .b(new_n12), .O(new_n54));
  nor2 g044(.a(new_n54), .b(new_n51), .O(new_n55));
  nor2 g045(.a(new_n55), .b(new_n48), .O(new_n56));
  nor2 g046(.a(_3), .b(new_n19), .O(new_n57));
  nor2 g047(.a(new_n15), .b(_9), .O(new_n58));
  nor2 g048(.a(new_n58), .b(new_n57), .O(new_n59));
  nor2 g049(.a(new_n13), .b(_8), .O(new_n60));
  inv1 g050(.a(new_n60), .O(new_n61));
  nor2 g051(.a(new_n61), .b(new_n20), .O(new_n62));
  inv1 g052(.a(new_n62), .O(new_n63));
  nor2 g053(.a(new_n63), .b(new_n59), .O(new_n64));
  nor2 g054(.a(new_n64), .b(new_n56), .O(new_n65));
  inv1 g055(.a(new_n65), .O(new_n66));
  nor2 g056(.a(new_n66), .b(new_n47), .O(new_n67));
  nor2 g057(.a(new_n67), .b(_1), .O(new_n68));
  inv1 g058(.a(_1), .O(new_n69));
  nor2 g059(.a(new_n12), .b(_8), .O(new_n70));
  nor2 g060(.a(_7), .b(new_n11), .O(new_n71));
  nor2 g061(.a(new_n71), .b(new_n70), .O(new_n72));
  inv1 g062(.a(new_n72), .O(new_n73));
  nor2 g063(.a(_4), .b(new_n19), .O(new_n74));
  nor2 g064(.a(new_n20), .b(_5), .O(new_n75));
  nor2 g065(.a(new_n75), .b(new_n74), .O(new_n76));
  inv1 g066(.a(new_n76), .O(new_n77));
  nor2 g067(.a(new_n77), .b(new_n73), .O(new_n78));
  nor2 g068(.a(new_n78), .b(new_n34), .O(new_n79));
  nor2 g069(.a(new_n61), .b(new_n50), .O(new_n80));
  nor2 g070(.a(new_n19), .b(_6), .O(new_n81));
  nor2 g071(.a(new_n81), .b(new_n75), .O(new_n82));
  nor2 g072(.a(new_n82), .b(new_n72), .O(new_n83));
  nor2 g073(.a(new_n83), .b(new_n80), .O(new_n84));
  inv1 g074(.a(new_n84), .O(new_n85));
  nor2 g075(.a(new_n85), .b(new_n79), .O(new_n86));
  nor2 g076(.a(new_n86), .b(new_n69), .O(new_n87));
  nor2 g077(.a(new_n69), .b(_3), .O(new_n88));
  nor2 g078(.a(_1), .b(new_n32), .O(new_n89));
  nor2 g079(.a(new_n89), .b(new_n58), .O(new_n90));
  inv1 g080(.a(new_n90), .O(new_n91));
  nor2 g081(.a(new_n91), .b(new_n88), .O(new_n92));
  inv1 g082(.a(new_n81), .O(new_n93));
  nor2 g083(.a(new_n93), .b(new_n20), .O(new_n94));
  inv1 g084(.a(new_n94), .O(new_n95));
  nor2 g085(.a(new_n95), .b(new_n92), .O(new_n96));
  nor2 g086(.a(_1), .b(new_n20), .O(new_n97));
  nor2 g087(.a(new_n69), .b(_4), .O(new_n98));
  nor2 g088(.a(new_n98), .b(new_n97), .O(new_n99));
  nor2 g089(.a(new_n48), .b(new_n13), .O(new_n100));
  inv1 g090(.a(new_n100), .O(new_n101));
  nor2 g091(.a(new_n101), .b(new_n99), .O(new_n102));
  nor2 g092(.a(new_n102), .b(new_n96), .O(new_n103));
  inv1 g093(.a(new_n103), .O(new_n104));
  nor2 g094(.a(new_n104), .b(new_n87), .O(new_n105));
  nor2 g095(.a(new_n105), .b(_2), .O(new_n106));
  nor2 g096(.a(new_n76), .b(_6), .O(new_n107));
  inv1 g097(.a(new_n107), .O(new_n108));
  nor2 g098(.a(_2), .b(new_n15), .O(new_n109));
  nor2 g099(.a(new_n49), .b(_3), .O(new_n110));
  nor2 g100(.a(new_n110), .b(new_n109), .O(new_n111));
  nor2 g101(.a(new_n111), .b(new_n69), .O(new_n112));
  inv1 g102(.a(new_n112), .O(new_n113));
  nor2 g103(.a(new_n113), .b(new_n108), .O(new_n114));
  nor2 g104(.a(new_n114), .b(new_n106), .O(new_n115));
  inv1 g105(.a(new_n115), .O(new_n116));
  nor2 g106(.a(new_n82), .b(new_n15), .O(new_n117));
  nor2 g107(.a(_1), .b(new_n19), .O(new_n118));
  inv1 g108(.a(new_n118), .O(new_n119));
  nor2 g109(.a(new_n119), .b(new_n13), .O(new_n120));
  nor2 g110(.a(new_n21), .b(new_n16), .O(new_n121));
  nor2 g111(.a(new_n121), .b(new_n49), .O(new_n122));
  nor2 g112(.a(new_n122), .b(new_n120), .O(new_n123));
  inv1 g113(.a(new_n123), .O(new_n124));
  nor2 g114(.a(new_n124), .b(new_n117), .O(new_n125));
  nor2 g115(.a(_7), .b(_8), .O(new_n126));
  inv1 g116(.a(new_n126), .O(new_n127));
  nor2 g117(.a(new_n127), .b(new_n125), .O(new_n128));
  inv1 g118(.a(new_n14), .O(new_n129));
  nor2 g119(.a(new_n129), .b(_1), .O(new_n130));
  nor2 g120(.a(new_n130), .b(new_n107), .O(new_n131));
  nor2 g121(.a(new_n131), .b(new_n72), .O(new_n132));
  nor2 g122(.a(_3), .b(_7), .O(new_n133));
  inv1 g123(.a(new_n133), .O(new_n134));
  nor2 g124(.a(new_n134), .b(new_n99), .O(new_n135));
  inv1 g125(.a(new_n16), .O(new_n136));
  nor2 g126(.a(_5), .b(new_n11), .O(new_n137));
  nor2 g127(.a(new_n137), .b(new_n74), .O(new_n138));
  inv1 g128(.a(new_n138), .O(new_n139));
  nor2 g129(.a(new_n139), .b(new_n136), .O(new_n140));
  nor2 g130(.a(new_n140), .b(new_n135), .O(new_n141));
  nor2 g131(.a(new_n141), .b(new_n13), .O(new_n142));
  nor2 g132(.a(new_n142), .b(new_n132), .O(new_n143));
  inv1 g133(.a(new_n143), .O(new_n144));
  nor2 g134(.a(new_n144), .b(new_n128), .O(new_n145));
  nor2 g135(.a(new_n145), .b(new_n32), .O(new_n146));
  nor2 g136(.a(_4), .b(new_n11), .O(new_n147));
  nor2 g137(.a(new_n147), .b(new_n97), .O(new_n148));
  nor2 g138(.a(_6), .b(new_n12), .O(new_n149));
  inv1 g139(.a(new_n149), .O(new_n150));
  nor2 g140(.a(new_n150), .b(new_n148), .O(new_n151));
  nor2 g141(.a(new_n72), .b(new_n129), .O(new_n152));
  nor2 g142(.a(new_n49), .b(_8), .O(new_n153));
  inv1 g143(.a(new_n153), .O(new_n154));
  nor2 g144(.a(new_n20), .b(_6), .O(new_n155));
  nor2 g145(.a(_3), .b(new_n13), .O(new_n156));
  nor2 g146(.a(new_n156), .b(new_n155), .O(new_n157));
  nor2 g147(.a(new_n157), .b(new_n154), .O(new_n158));
  nor2 g148(.a(new_n158), .b(new_n152), .O(new_n159));
  inv1 g149(.a(new_n159), .O(new_n160));
  nor2 g150(.a(new_n160), .b(new_n151), .O(new_n161));
  nor2 g151(.a(new_n161), .b(new_n19), .O(new_n162));
  nor2 g152(.a(new_n138), .b(_2), .O(new_n163));
  nor2 g153(.a(new_n36), .b(_3), .O(new_n164));
  nor2 g154(.a(_5), .b(_7), .O(new_n165));
  inv1 g155(.a(new_n165), .O(new_n166));
  nor2 g156(.a(new_n166), .b(new_n49), .O(new_n167));
  nor2 g157(.a(new_n167), .b(new_n164), .O(new_n168));
  inv1 g158(.a(new_n168), .O(new_n169));
  nor2 g159(.a(new_n169), .b(new_n163), .O(new_n170));
  nor2 g160(.a(new_n69), .b(new_n13), .O(new_n171));
  inv1 g161(.a(new_n171), .O(new_n172));
  nor2 g162(.a(new_n172), .b(new_n170), .O(new_n173));
  nor2 g163(.a(new_n154), .b(new_n69), .O(new_n174));
  inv1 g164(.a(new_n155), .O(new_n175));
  nor2 g165(.a(new_n175), .b(new_n11), .O(new_n176));
  nor2 g166(.a(new_n176), .b(new_n174), .O(new_n177));
  nor2 g167(.a(new_n15), .b(_7), .O(new_n178));
  inv1 g168(.a(new_n178), .O(new_n179));
  nor2 g169(.a(new_n179), .b(new_n177), .O(new_n180));
  nor2 g170(.a(_2), .b(new_n11), .O(new_n181));
  nor2 g171(.a(new_n60), .b(new_n41), .O(new_n182));
  inv1 g172(.a(new_n182), .O(new_n183));
  nor2 g173(.a(new_n183), .b(new_n181), .O(new_n184));
  nor2 g174(.a(_5), .b(new_n12), .O(new_n185));
  inv1 g175(.a(new_n185), .O(new_n186));
  nor2 g176(.a(new_n186), .b(new_n20), .O(new_n187));
  inv1 g177(.a(new_n187), .O(new_n188));
  nor2 g178(.a(new_n188), .b(new_n184), .O(new_n189));
  nor2 g179(.a(new_n189), .b(new_n180), .O(new_n190));
  inv1 g180(.a(new_n190), .O(new_n191));
  nor2 g181(.a(new_n191), .b(new_n173), .O(new_n192));
  inv1 g182(.a(new_n192), .O(new_n193));
  nor2 g183(.a(new_n193), .b(new_n162), .O(new_n194));
  nor2 g184(.a(new_n194), .b(_9), .O(new_n195));
  nor2 g185(.a(new_n195), .b(new_n146), .O(new_n196));
  inv1 g186(.a(new_n196), .O(new_n197));
  nor2 g187(.a(new_n197), .b(new_n116), .O(new_n198));
  inv1 g188(.a(new_n198), .O(new_n199));
  nor2 g189(.a(new_n70), .b(new_n38), .O(new_n200));
  nor2 g190(.a(new_n200), .b(new_n34), .O(new_n201));
  nor2 g191(.a(new_n15), .b(new_n11), .O(new_n202));
  inv1 g192(.a(new_n97), .O(new_n203));
  nor2 g193(.a(new_n133), .b(new_n203), .O(new_n204));
  inv1 g194(.a(new_n204), .O(new_n205));
  nor2 g195(.a(new_n205), .b(new_n202), .O(new_n206));
  inv1 g196(.a(new_n98), .O(new_n207));
  nor2 g197(.a(new_n186), .b(new_n207), .O(new_n208));
  nor2 g198(.a(new_n208), .b(new_n206), .O(new_n209));
  inv1 g199(.a(new_n209), .O(new_n210));
  nor2 g200(.a(new_n210), .b(new_n201), .O(new_n211));
  nor2 g201(.a(new_n211), .b(_6), .O(new_n212));
  nor2 g202(.a(new_n155), .b(new_n38), .O(new_n213));
  inv1 g203(.a(new_n213), .O(new_n214));
  nor2 g204(.a(new_n214), .b(new_n185), .O(new_n215));
  nor2 g205(.a(new_n11), .b(_9), .O(new_n216));
  inv1 g206(.a(new_n216), .O(new_n217));
  nor2 g207(.a(new_n217), .b(new_n215), .O(new_n218));
  nor2 g208(.a(new_n71), .b(new_n52), .O(new_n219));
  nor2 g209(.a(_5), .b(new_n13), .O(new_n220));
  inv1 g210(.a(new_n220), .O(new_n221));
  nor2 g211(.a(new_n221), .b(new_n219), .O(new_n222));
  nor2 g212(.a(new_n69), .b(_5), .O(new_n223));
  nor2 g213(.a(_1), .b(new_n11), .O(new_n224));
  nor2 g214(.a(new_n224), .b(new_n223), .O(new_n225));
  nor2 g215(.a(_4), .b(new_n32), .O(new_n226));
  inv1 g216(.a(new_n226), .O(new_n227));
  nor2 g217(.a(new_n227), .b(new_n225), .O(new_n228));
  nor2 g218(.a(new_n228), .b(new_n222), .O(new_n229));
  inv1 g219(.a(new_n229), .O(new_n230));
  nor2 g220(.a(new_n230), .b(new_n218), .O(new_n231));
  nor2 g221(.a(new_n231), .b(_3), .O(new_n232));
  nor2 g222(.a(new_n221), .b(_1), .O(new_n233));
  inv1 g223(.a(new_n233), .O(new_n234));
  nor2 g224(.a(new_n234), .b(new_n121), .O(new_n235));
  nor2 g225(.a(new_n235), .b(new_n232), .O(new_n236));
  inv1 g226(.a(new_n236), .O(new_n237));
  nor2 g227(.a(new_n237), .b(new_n212), .O(new_n238));
  nor2 g228(.a(new_n238), .b(new_n49), .O(new_n239));
  nor2 g229(.a(new_n110), .b(new_n24), .O(new_n240));
  nor2 g230(.a(new_n13), .b(_9), .O(new_n241));
  inv1 g231(.a(new_n241), .O(new_n242));
  nor2 g232(.a(new_n242), .b(new_n240), .O(new_n243));
  inv1 g233(.a(new_n109), .O(new_n244));
  nor2 g234(.a(new_n225), .b(new_n244), .O(new_n245));
  inv1 g235(.a(new_n57), .O(new_n246));
  nor2 g236(.a(new_n154), .b(new_n246), .O(new_n247));
  nor2 g237(.a(new_n247), .b(new_n245), .O(new_n248));
  inv1 g238(.a(new_n248), .O(new_n249));
  nor2 g239(.a(new_n249), .b(new_n243), .O(new_n250));
  nor2 g240(.a(new_n250), .b(new_n12), .O(new_n251));
  nor2 g241(.a(new_n13), .b(_7), .O(new_n252));
  nor2 g242(.a(new_n49), .b(_6), .O(new_n253));
  nor2 g243(.a(new_n253), .b(new_n70), .O(new_n254));
  inv1 g244(.a(new_n254), .O(new_n255));
  nor2 g245(.a(new_n255), .b(new_n252), .O(new_n256));
  nor2 g246(.a(new_n256), .b(new_n119), .O(new_n257));
  nor2 g247(.a(new_n69), .b(_2), .O(new_n258));
  inv1 g248(.a(new_n258), .O(new_n259));
  nor2 g249(.a(new_n259), .b(new_n219), .O(new_n260));
  nor2 g250(.a(new_n49), .b(_9), .O(new_n261));
  inv1 g251(.a(new_n261), .O(new_n262));
  nor2 g252(.a(new_n262), .b(new_n72), .O(new_n263));
  nor2 g253(.a(new_n263), .b(new_n260), .O(new_n264));
  inv1 g254(.a(new_n264), .O(new_n265));
  nor2 g255(.a(new_n265), .b(new_n257), .O(new_n266));
  nor2 g256(.a(new_n266), .b(new_n15), .O(new_n267));
  nor2 g257(.a(new_n69), .b(new_n11), .O(new_n268));
  inv1 g258(.a(new_n268), .O(new_n269));
  nor2 g259(.a(new_n269), .b(new_n168), .O(new_n270));
  nor2 g260(.a(new_n270), .b(new_n267), .O(new_n271));
  inv1 g261(.a(new_n271), .O(new_n272));
  nor2 g262(.a(new_n272), .b(new_n251), .O(new_n273));
  nor2 g263(.a(new_n273), .b(_4), .O(new_n274));
  nor2 g264(.a(new_n274), .b(new_n239), .O(new_n275));
  inv1 g265(.a(new_n275), .O(new_n276));
  nor2 g266(.a(new_n276), .b(new_n199), .O(new_n277));
  inv1 g267(.a(new_n277), .O(new_n278));
  nor2 g268(.a(new_n278), .b(new_n68), .O(new_n279));
  inv1 g269(.a(new_n279), .O(_52));
endmodule


